`timescale 1ns / 1ps
module supra2(
input enable,
input clock,
input [9:0] posx, posy,
input [9:0] hcount,
input [9:0] vcount,
output reg[2:0] red,
output reg[2:0] green,
output reg[1:0] blue,
output reg data);

always @(posedge clock)
begin
	if(enable)
	begin
		if(hcount >= posx & hcount < posx + RESOLUCION_X & vcount >= posy & vcount < posy + RESOLUCION_Y)
		begin
			if (supra2[vcount - posy][hcount - posx][8] == 1'b1)
			begin
				red   <= supra2[vcount- posy][hcount- posx][7:5];
				green <= supra2[vcount- posy][hcount- posx][4:2];
            blue 	<= supra2[vcount- posy][hcount- posx][1:0];
				data  <= 1'b1;
			end
			else
				data <= 0;
			end
		else
		data <= 0;
	end
end

parameter RESOLUCION_X = 18;
parameter RESOLUCION_Y = 45;
wire [8:0] supra2[RESOLUCION_Y - 1'b1 : 0][RESOLUCION_X - 1'b1 : 0];
assign supra2[0][4] = 9'b111101000;
assign supra2[0][5] = 9'b111101000;
assign supra2[0][6] = 9'b111101000;
assign supra2[0][7] = 9'b111101000;
assign supra2[0][8] = 9'b111101000;
assign supra2[0][9] = 9'b111101000;
assign supra2[0][10] = 9'b111101000;
assign supra2[0][11] = 9'b111101000;
assign supra2[0][12] = 9'b111101000;
assign supra2[0][13] = 9'b111101000;
assign supra2[1][3] = 9'b111101000;
assign supra2[1][4] = 9'b110110001;
assign supra2[1][5] = 9'b110010110;
assign supra2[1][6] = 9'b111101000;
assign supra2[1][7] = 9'b111101000;
assign supra2[1][8] = 9'b111101000;
assign supra2[1][9] = 9'b111101000;
assign supra2[1][10] = 9'b111101000;
assign supra2[1][11] = 9'b111101000;
assign supra2[1][12] = 9'b110010110;
assign supra2[1][13] = 9'b110110001;
assign supra2[1][14] = 9'b111101000;
assign supra2[2][2] = 9'b111101000;
assign supra2[2][3] = 9'b110010110;
assign supra2[2][4] = 9'b101111111;
assign supra2[2][5] = 9'b110010110;
assign supra2[2][6] = 9'b111101000;
assign supra2[2][7] = 9'b111101000;
assign supra2[2][8] = 9'b111101000;
assign supra2[2][9] = 9'b111101000;
assign supra2[2][10] = 9'b111101000;
assign supra2[2][11] = 9'b111101000;
assign supra2[2][12] = 9'b110010010;
assign supra2[2][13] = 9'b101111111;
assign supra2[2][14] = 9'b110010110;
assign supra2[2][15] = 9'b111101000;
assign supra2[3][1] = 9'b111100100;
assign supra2[3][2] = 9'b110110001;
assign supra2[3][3] = 9'b101110111;
assign supra2[3][4] = 9'b110101101;
assign supra2[3][5] = 9'b111101000;
assign supra2[3][6] = 9'b111101000;
assign supra2[3][7] = 9'b111101000;
assign supra2[3][8] = 9'b111101000;
assign supra2[3][9] = 9'b111101000;
assign supra2[3][10] = 9'b111101000;
assign supra2[3][11] = 9'b111101000;
assign supra2[3][12] = 9'b111101000;
assign supra2[3][13] = 9'b110101101;
assign supra2[3][14] = 9'b101110111;
assign supra2[3][15] = 9'b110110001;
assign supra2[3][16] = 9'b111100100;
assign supra2[4][1] = 9'b111101000;
assign supra2[4][2] = 9'b111101100;
assign supra2[4][3] = 9'b111101000;
assign supra2[4][4] = 9'b111101000;
assign supra2[4][5] = 9'b111101000;
assign supra2[4][6] = 9'b111101000;
assign supra2[4][7] = 9'b111101000;
assign supra2[4][8] = 9'b111101000;
assign supra2[4][9] = 9'b111101000;
assign supra2[4][10] = 9'b111101000;
assign supra2[4][11] = 9'b111101000;
assign supra2[4][12] = 9'b111101000;
assign supra2[4][13] = 9'b111101000;
assign supra2[4][14] = 9'b111101000;
assign supra2[4][15] = 9'b111101000;
assign supra2[4][16] = 9'b111101000;
assign supra2[5][1] = 9'b111101000;
assign supra2[5][2] = 9'b111101000;
assign supra2[5][3] = 9'b111101000;
assign supra2[5][4] = 9'b111101000;
assign supra2[5][5] = 9'b111101000;
assign supra2[5][6] = 9'b111101000;
assign supra2[5][7] = 9'b111101000;
assign supra2[5][8] = 9'b111101000;
assign supra2[5][9] = 9'b111101000;
assign supra2[5][10] = 9'b111101000;
assign supra2[5][11] = 9'b111101000;
assign supra2[5][12] = 9'b111101000;
assign supra2[5][13] = 9'b111101000;
assign supra2[5][14] = 9'b111101000;
assign supra2[5][15] = 9'b111101000;
assign supra2[5][16] = 9'b111101000;
assign supra2[6][1] = 9'b111101000;
assign supra2[6][2] = 9'b111101000;
assign supra2[6][3] = 9'b111101000;
assign supra2[6][4] = 9'b111101000;
assign supra2[6][5] = 9'b111101000;
assign supra2[6][6] = 9'b111101000;
assign supra2[6][7] = 9'b111101000;
assign supra2[6][8] = 9'b111101000;
assign supra2[6][9] = 9'b111101000;
assign supra2[6][10] = 9'b111101000;
assign supra2[6][11] = 9'b111101000;
assign supra2[6][12] = 9'b111101000;
assign supra2[6][13] = 9'b111101000;
assign supra2[6][14] = 9'b111101000;
assign supra2[6][15] = 9'b111101000;
assign supra2[6][16] = 9'b111101000;
assign supra2[7][1] = 9'b111101000;
assign supra2[7][2] = 9'b111101000;
assign supra2[7][3] = 9'b111101000;
assign supra2[7][4] = 9'b111101000;
assign supra2[7][5] = 9'b111101000;
assign supra2[7][6] = 9'b111101000;
assign supra2[7][7] = 9'b111101000;
assign supra2[7][8] = 9'b111101000;
assign supra2[7][9] = 9'b111101000;
assign supra2[7][10] = 9'b111101000;
assign supra2[7][11] = 9'b111101000;
assign supra2[7][12] = 9'b111101000;
assign supra2[7][13] = 9'b111101000;
assign supra2[7][14] = 9'b111101000;
assign supra2[7][15] = 9'b111101000;
assign supra2[7][16] = 9'b111101000;
assign supra2[8][1] = 9'b111101000;
assign supra2[8][2] = 9'b111101000;
assign supra2[8][3] = 9'b111101000;
assign supra2[8][4] = 9'b111101000;
assign supra2[8][5] = 9'b111101000;
assign supra2[8][6] = 9'b111101000;
assign supra2[8][7] = 9'b111101000;
assign supra2[8][8] = 9'b111101000;
assign supra2[8][9] = 9'b111101000;
assign supra2[8][10] = 9'b111101000;
assign supra2[8][11] = 9'b111101000;
assign supra2[8][12] = 9'b111101000;
assign supra2[8][13] = 9'b111101000;
assign supra2[8][14] = 9'b111101000;
assign supra2[8][15] = 9'b111101000;
assign supra2[8][16] = 9'b111101000;
assign supra2[9][1] = 9'b111101000;
assign supra2[9][2] = 9'b111101000;
assign supra2[9][3] = 9'b111101000;
assign supra2[9][4] = 9'b111101000;
assign supra2[9][5] = 9'b111101000;
assign supra2[9][6] = 9'b111101000;
assign supra2[9][7] = 9'b111101000;
assign supra2[9][8] = 9'b111101000;
assign supra2[9][9] = 9'b111101000;
assign supra2[9][10] = 9'b111101000;
assign supra2[9][11] = 9'b111101000;
assign supra2[9][12] = 9'b111101000;
assign supra2[9][13] = 9'b111101000;
assign supra2[9][14] = 9'b111101000;
assign supra2[9][15] = 9'b111101000;
assign supra2[9][16] = 9'b111101000;
assign supra2[10][1] = 9'b111101000;
assign supra2[10][2] = 9'b111101000;
assign supra2[10][3] = 9'b111101000;
assign supra2[10][4] = 9'b111101000;
assign supra2[10][5] = 9'b111101000;
assign supra2[10][6] = 9'b111101000;
assign supra2[10][7] = 9'b111101000;
assign supra2[10][8] = 9'b111101000;
assign supra2[10][9] = 9'b111101000;
assign supra2[10][10] = 9'b111101000;
assign supra2[10][11] = 9'b111101000;
assign supra2[10][12] = 9'b111101000;
assign supra2[10][13] = 9'b111101000;
assign supra2[10][14] = 9'b111101000;
assign supra2[10][15] = 9'b111101000;
assign supra2[10][16] = 9'b111101000;
assign supra2[10][17] = 9'b111101000;
assign supra2[11][0] = 9'b111101000;
assign supra2[11][1] = 9'b111101000;
assign supra2[11][2] = 9'b111101000;
assign supra2[11][3] = 9'b111101000;
assign supra2[11][4] = 9'b111101000;
assign supra2[11][5] = 9'b111101000;
assign supra2[11][6] = 9'b111101000;
assign supra2[11][7] = 9'b111101000;
assign supra2[11][8] = 9'b111101000;
assign supra2[11][9] = 9'b111101000;
assign supra2[11][10] = 9'b111101000;
assign supra2[11][11] = 9'b111101000;
assign supra2[11][12] = 9'b111101000;
assign supra2[11][13] = 9'b111101000;
assign supra2[11][14] = 9'b111101000;
assign supra2[11][15] = 9'b111101000;
assign supra2[11][16] = 9'b111101000;
assign supra2[11][17] = 9'b111101000;
assign supra2[12][0] = 9'b111101000;
assign supra2[12][1] = 9'b111101000;
assign supra2[12][2] = 9'b111101000;
assign supra2[12][3] = 9'b111101000;
assign supra2[12][4] = 9'b111101000;
assign supra2[12][5] = 9'b111101000;
assign supra2[12][6] = 9'b111101000;
assign supra2[12][7] = 9'b111101000;
assign supra2[12][8] = 9'b111101000;
assign supra2[12][9] = 9'b111101000;
assign supra2[12][10] = 9'b111101000;
assign supra2[12][11] = 9'b111101000;
assign supra2[12][12] = 9'b111101000;
assign supra2[12][13] = 9'b111101000;
assign supra2[12][14] = 9'b111101000;
assign supra2[12][15] = 9'b111101000;
assign supra2[12][16] = 9'b111101000;
assign supra2[12][17] = 9'b111101000;
assign supra2[13][0] = 9'b111101000;
assign supra2[13][1] = 9'b111101000;
assign supra2[13][2] = 9'b111101000;
assign supra2[13][3] = 9'b111101000;
assign supra2[13][4] = 9'b111101000;
assign supra2[13][5] = 9'b111101000;
assign supra2[13][6] = 9'b111101000;
assign supra2[13][7] = 9'b110101000;
assign supra2[13][8] = 9'b110101000;
assign supra2[13][9] = 9'b110101000;
assign supra2[13][10] = 9'b110101000;
assign supra2[13][11] = 9'b111101000;
assign supra2[13][12] = 9'b111101000;
assign supra2[13][13] = 9'b111101000;
assign supra2[13][14] = 9'b111101000;
assign supra2[13][15] = 9'b111101000;
assign supra2[13][16] = 9'b111101000;
assign supra2[13][17] = 9'b111101000;
assign supra2[14][0] = 9'b111101000;
assign supra2[14][1] = 9'b111101000;
assign supra2[14][2] = 9'b111101000;
assign supra2[14][3] = 9'b111101000;
assign supra2[14][4] = 9'b101100100;
assign supra2[14][5] = 9'b101000100;
assign supra2[14][6] = 9'b100100000;
assign supra2[14][7] = 9'b100000000;
assign supra2[14][8] = 9'b100000000;
assign supra2[14][9] = 9'b100000000;
assign supra2[14][10] = 9'b100000000;
assign supra2[14][11] = 9'b100100000;
assign supra2[14][12] = 9'b101000100;
assign supra2[14][13] = 9'b101100100;
assign supra2[14][14] = 9'b111101000;
assign supra2[14][15] = 9'b111101000;
assign supra2[14][16] = 9'b111101000;
assign supra2[14][17] = 9'b111101000;
assign supra2[15][0] = 9'b111101000;
assign supra2[15][1] = 9'b111101000;
assign supra2[15][2] = 9'b111101000;
assign supra2[15][3] = 9'b100100000;
assign supra2[15][4] = 9'b100000000;
assign supra2[15][5] = 9'b100000000;
assign supra2[15][6] = 9'b100000100;
assign supra2[15][7] = 9'b100000101;
assign supra2[15][8] = 9'b100000101;
assign supra2[15][9] = 9'b100000101;
assign supra2[15][10] = 9'b100000101;
assign supra2[15][11] = 9'b100000100;
assign supra2[15][12] = 9'b100000000;
assign supra2[15][13] = 9'b100000000;
assign supra2[15][14] = 9'b100100000;
assign supra2[15][15] = 9'b111101000;
assign supra2[15][16] = 9'b111101000;
assign supra2[15][17] = 9'b111101000;
assign supra2[16][1] = 9'b111101000;
assign supra2[16][2] = 9'b101000100;
assign supra2[16][3] = 9'b100000100;
assign supra2[16][4] = 9'b100001001;
assign supra2[16][5] = 9'b100001010;
assign supra2[16][6] = 9'b100001111;
assign supra2[16][7] = 9'b100001111;
assign supra2[16][8] = 9'b100001111;
assign supra2[16][9] = 9'b100001111;
assign supra2[16][10] = 9'b100001111;
assign supra2[16][11] = 9'b100001111;
assign supra2[16][12] = 9'b100001111;
assign supra2[16][13] = 9'b100001011;
assign supra2[16][14] = 9'b100000101;
assign supra2[16][15] = 9'b101000100;
assign supra2[16][16] = 9'b111101000;
assign supra2[17][1] = 9'b111101000;
assign supra2[17][2] = 9'b101001000;
assign supra2[17][3] = 9'b100001111;
assign supra2[17][4] = 9'b100001111;
assign supra2[17][5] = 9'b100001111;
assign supra2[17][6] = 9'b100001111;
assign supra2[17][7] = 9'b100001111;
assign supra2[17][8] = 9'b100001111;
assign supra2[17][9] = 9'b100001111;
assign supra2[17][10] = 9'b100001111;
assign supra2[17][11] = 9'b100001111;
assign supra2[17][12] = 9'b100001111;
assign supra2[17][13] = 9'b100001111;
assign supra2[17][14] = 9'b100001111;
assign supra2[17][15] = 9'b101001000;
assign supra2[17][16] = 9'b111101000;
assign supra2[18][1] = 9'b111101000;
assign supra2[18][2] = 9'b101101000;
assign supra2[18][3] = 9'b100001111;
assign supra2[18][4] = 9'b100001111;
assign supra2[18][5] = 9'b100001111;
assign supra2[18][6] = 9'b100001111;
assign supra2[18][7] = 9'b100001111;
assign supra2[18][8] = 9'b100001111;
assign supra2[18][9] = 9'b100001111;
assign supra2[18][10] = 9'b100001111;
assign supra2[18][11] = 9'b100001111;
assign supra2[18][12] = 9'b100001111;
assign supra2[18][13] = 9'b100001111;
assign supra2[18][14] = 9'b100001111;
assign supra2[18][15] = 9'b101101000;
assign supra2[18][16] = 9'b111101000;
assign supra2[19][0] = 9'b111101000;
assign supra2[19][1] = 9'b111101000;
assign supra2[19][2] = 9'b101101001;
assign supra2[19][3] = 9'b100000101;
assign supra2[19][4] = 9'b100000110;
assign supra2[19][5] = 9'b100001111;
assign supra2[19][6] = 9'b100001011;
assign supra2[19][7] = 9'b100000110;
assign supra2[19][8] = 9'b100001011;
assign supra2[19][9] = 9'b100001111;
assign supra2[19][10] = 9'b100000110;
assign supra2[19][11] = 9'b100000001;
assign supra2[19][12] = 9'b100000001;
assign supra2[19][13] = 9'b100000001;
assign supra2[19][14] = 9'b100000101;
assign supra2[19][15] = 9'b101101001;
assign supra2[19][16] = 9'b111101000;
assign supra2[19][17] = 9'b111101000;
assign supra2[20][0] = 9'b111101000;
assign supra2[20][1] = 9'b111101000;
assign supra2[20][2] = 9'b101001101;
assign supra2[20][3] = 9'b100100100;
assign supra2[20][4] = 9'b100000110;
assign supra2[20][5] = 9'b100001011;
assign supra2[20][6] = 9'b100000101;
assign supra2[20][7] = 9'b100000001;
assign supra2[20][8] = 9'b100001111;
assign supra2[20][9] = 9'b100001111;
assign supra2[20][10] = 9'b100000101;
assign supra2[20][11] = 9'b100000110;
assign supra2[20][12] = 9'b100000110;
assign supra2[20][13] = 9'b100000111;
assign supra2[20][14] = 9'b100100101;
assign supra2[20][15] = 9'b101001001;
assign supra2[20][16] = 9'b111101000;
assign supra2[20][17] = 9'b111101000;
assign supra2[21][1] = 9'b111101000;
assign supra2[21][2] = 9'b100001010;
assign supra2[21][3] = 9'b101001001;
assign supra2[21][4] = 9'b100001111;
assign supra2[21][5] = 9'b100001111;
assign supra2[21][6] = 9'b100001111;
assign supra2[21][7] = 9'b100001010;
assign supra2[21][8] = 9'b100001011;
assign supra2[21][9] = 9'b100001011;
assign supra2[21][10] = 9'b100001010;
assign supra2[21][11] = 9'b100001111;
assign supra2[21][12] = 9'b100001111;
assign supra2[21][13] = 9'b100001111;
assign supra2[21][14] = 9'b101001001;
assign supra2[21][15] = 9'b100001010;
assign supra2[21][16] = 9'b111101000;
assign supra2[22][1] = 9'b111101000;
assign supra2[22][2] = 9'b100001111;
assign supra2[22][3] = 9'b101101001;
assign supra2[22][4] = 9'b110101000;
assign supra2[22][5] = 9'b110001000;
assign supra2[22][6] = 9'b110101000;
assign supra2[22][7] = 9'b110101000;
assign supra2[22][8] = 9'b111101000;
assign supra2[22][9] = 9'b111101000;
assign supra2[22][10] = 9'b110101000;
assign supra2[22][11] = 9'b110101000;
assign supra2[22][12] = 9'b110001000;
assign supra2[22][13] = 9'b110101000;
assign supra2[22][14] = 9'b101101001;
assign supra2[22][15] = 9'b100001111;
assign supra2[22][16] = 9'b111101000;
assign supra2[23][1] = 9'b111101000;
assign supra2[23][2] = 9'b100001111;
assign supra2[23][3] = 9'b100101110;
assign supra2[23][4] = 9'b111101000;
assign supra2[23][5] = 9'b111101000;
assign supra2[23][6] = 9'b111101000;
assign supra2[23][7] = 9'b111101000;
assign supra2[23][8] = 9'b111101000;
assign supra2[23][9] = 9'b111101000;
assign supra2[23][10] = 9'b111101000;
assign supra2[23][11] = 9'b111101000;
assign supra2[23][12] = 9'b111101000;
assign supra2[23][13] = 9'b111101000;
assign supra2[23][14] = 9'b100101110;
assign supra2[23][15] = 9'b100001111;
assign supra2[23][16] = 9'b111101000;
assign supra2[24][1] = 9'b111101000;
assign supra2[24][2] = 9'b100001011;
assign supra2[24][3] = 9'b100001110;
assign supra2[24][4] = 9'b111101000;
assign supra2[24][5] = 9'b111101000;
assign supra2[24][6] = 9'b111101000;
assign supra2[24][7] = 9'b111101000;
assign supra2[24][8] = 9'b111101000;
assign supra2[24][9] = 9'b111101000;
assign supra2[24][10] = 9'b111101000;
assign supra2[24][11] = 9'b111101000;
assign supra2[24][12] = 9'b111101000;
assign supra2[24][13] = 9'b111101000;
assign supra2[24][14] = 9'b100101110;
assign supra2[24][15] = 9'b100001011;
assign supra2[24][16] = 9'b111101000;
assign supra2[25][1] = 9'b111101000;
assign supra2[25][2] = 9'b100001111;
assign supra2[25][3] = 9'b100001111;
assign supra2[25][4] = 9'b111101000;
assign supra2[25][5] = 9'b111101000;
assign supra2[25][6] = 9'b111101000;
assign supra2[25][7] = 9'b111101000;
assign supra2[25][8] = 9'b111101000;
assign supra2[25][9] = 9'b111101000;
assign supra2[25][10] = 9'b111101000;
assign supra2[25][11] = 9'b111101000;
assign supra2[25][12] = 9'b111101000;
assign supra2[25][13] = 9'b111101000;
assign supra2[25][14] = 9'b100001111;
assign supra2[25][15] = 9'b100001111;
assign supra2[25][16] = 9'b111101000;
assign supra2[26][1] = 9'b111101000;
assign supra2[26][2] = 9'b100001111;
assign supra2[26][3] = 9'b100001111;
assign supra2[26][4] = 9'b111101000;
assign supra2[26][5] = 9'b111101000;
assign supra2[26][6] = 9'b111101000;
assign supra2[26][7] = 9'b111101000;
assign supra2[26][8] = 9'b111101000;
assign supra2[26][9] = 9'b111101000;
assign supra2[26][10] = 9'b111101000;
assign supra2[26][11] = 9'b111101000;
assign supra2[26][12] = 9'b111101000;
assign supra2[26][13] = 9'b111101000;
assign supra2[26][14] = 9'b100101111;
assign supra2[26][15] = 9'b100001111;
assign supra2[26][16] = 9'b111101000;
assign supra2[27][1] = 9'b111101000;
assign supra2[27][2] = 9'b100001010;
assign supra2[27][3] = 9'b100101010;
assign supra2[27][4] = 9'b111101000;
assign supra2[27][5] = 9'b111101000;
assign supra2[27][6] = 9'b111101000;
assign supra2[27][7] = 9'b111101000;
assign supra2[27][8] = 9'b111101000;
assign supra2[27][9] = 9'b111101000;
assign supra2[27][10] = 9'b111101000;
assign supra2[27][11] = 9'b111101000;
assign supra2[27][12] = 9'b111101000;
assign supra2[27][13] = 9'b111101000;
assign supra2[27][14] = 9'b100101010;
assign supra2[27][15] = 9'b100001010;
assign supra2[27][16] = 9'b111101000;
assign supra2[28][1] = 9'b111101000;
assign supra2[28][2] = 9'b100000101;
assign supra2[28][3] = 9'b100100101;
assign supra2[28][4] = 9'b111101000;
assign supra2[28][5] = 9'b111101000;
assign supra2[28][6] = 9'b111101000;
assign supra2[28][7] = 9'b111101000;
assign supra2[28][8] = 9'b111101000;
assign supra2[28][9] = 9'b111101000;
assign supra2[28][10] = 9'b111101000;
assign supra2[28][11] = 9'b111101000;
assign supra2[28][12] = 9'b111101000;
assign supra2[28][13] = 9'b111101000;
assign supra2[28][14] = 9'b101000101;
assign supra2[28][15] = 9'b100000101;
assign supra2[28][16] = 9'b111101000;
assign supra2[29][1] = 9'b111101000;
assign supra2[29][2] = 9'b100000101;
assign supra2[29][3] = 9'b101000100;
assign supra2[29][4] = 9'b111101000;
assign supra2[29][5] = 9'b111101000;
assign supra2[29][6] = 9'b111101000;
assign supra2[29][7] = 9'b111101000;
assign supra2[29][8] = 9'b111101000;
assign supra2[29][9] = 9'b111101000;
assign supra2[29][10] = 9'b111101000;
assign supra2[29][11] = 9'b111101000;
assign supra2[29][12] = 9'b111101000;
assign supra2[29][13] = 9'b111101000;
assign supra2[29][14] = 9'b101100100;
assign supra2[29][15] = 9'b100000101;
assign supra2[29][16] = 9'b111101000;
assign supra2[30][0] = 9'b111101000;
assign supra2[30][1] = 9'b111101000;
assign supra2[30][2] = 9'b100001010;
assign supra2[30][3] = 9'b110001000;
assign supra2[30][4] = 9'b111101000;
assign supra2[30][5] = 9'b111101000;
assign supra2[30][6] = 9'b111101000;
assign supra2[30][7] = 9'b111101000;
assign supra2[30][8] = 9'b111101000;
assign supra2[30][9] = 9'b111101000;
assign supra2[30][10] = 9'b111101000;
assign supra2[30][11] = 9'b111101000;
assign supra2[30][12] = 9'b111101000;
assign supra2[30][13] = 9'b111101000;
assign supra2[30][14] = 9'b110001000;
assign supra2[30][15] = 9'b100001010;
assign supra2[30][16] = 9'b111101000;
assign supra2[30][17] = 9'b111101000;
assign supra2[31][0] = 9'b111101000;
assign supra2[31][1] = 9'b111101000;
assign supra2[31][2] = 9'b101101001;
assign supra2[31][3] = 9'b111101000;
assign supra2[31][4] = 9'b110001000;
assign supra2[31][5] = 9'b101001000;
assign supra2[31][6] = 9'b101001000;
assign supra2[31][7] = 9'b101001000;
assign supra2[31][8] = 9'b101101000;
assign supra2[31][9] = 9'b101101000;
assign supra2[31][10] = 9'b101001000;
assign supra2[31][11] = 9'b101001000;
assign supra2[31][12] = 9'b101001000;
assign supra2[31][13] = 9'b110001000;
assign supra2[31][14] = 9'b111101000;
assign supra2[31][15] = 9'b101001001;
assign supra2[31][16] = 9'b111101000;
assign supra2[31][17] = 9'b111101000;
assign supra2[32][0] = 9'b111101000;
assign supra2[32][1] = 9'b111101000;
assign supra2[32][2] = 9'b111101000;
assign supra2[32][3] = 9'b111101000;
assign supra2[32][4] = 9'b100001001;
assign supra2[32][5] = 9'b100001111;
assign supra2[32][6] = 9'b100001111;
assign supra2[32][7] = 9'b100001111;
assign supra2[32][8] = 9'b100001111;
assign supra2[32][9] = 9'b100001111;
assign supra2[32][10] = 9'b100001111;
assign supra2[32][11] = 9'b100001111;
assign supra2[32][12] = 9'b100001111;
assign supra2[32][13] = 9'b100001001;
assign supra2[32][14] = 9'b111101000;
assign supra2[32][15] = 9'b111101000;
assign supra2[32][16] = 9'b111101000;
assign supra2[32][17] = 9'b111101000;
assign supra2[33][0] = 9'b111101000;
assign supra2[33][1] = 9'b111101000;
assign supra2[33][2] = 9'b111101000;
assign supra2[33][3] = 9'b110101000;
assign supra2[33][4] = 9'b100001111;
assign supra2[33][5] = 9'b100001111;
assign supra2[33][6] = 9'b100001111;
assign supra2[33][7] = 9'b100001111;
assign supra2[33][8] = 9'b100001111;
assign supra2[33][9] = 9'b100001111;
assign supra2[33][10] = 9'b100001111;
assign supra2[33][11] = 9'b100001111;
assign supra2[33][12] = 9'b100001111;
assign supra2[33][13] = 9'b100001111;
assign supra2[33][14] = 9'b110001000;
assign supra2[33][15] = 9'b111101000;
assign supra2[33][16] = 9'b111101000;
assign supra2[33][17] = 9'b111101000;
assign supra2[34][0] = 9'b111101000;
assign supra2[34][1] = 9'b111101000;
assign supra2[34][2] = 9'b111101000;
assign supra2[34][3] = 9'b110001000;
assign supra2[34][4] = 9'b100001111;
assign supra2[34][5] = 9'b100001111;
assign supra2[34][6] = 9'b100001111;
assign supra2[34][7] = 9'b100001111;
assign supra2[34][8] = 9'b100001111;
assign supra2[34][9] = 9'b100001111;
assign supra2[34][10] = 9'b100001111;
assign supra2[34][11] = 9'b100001111;
assign supra2[34][12] = 9'b100001111;
assign supra2[34][13] = 9'b100001111;
assign supra2[34][14] = 9'b110001000;
assign supra2[34][15] = 9'b111101000;
assign supra2[34][16] = 9'b111101000;
assign supra2[34][17] = 9'b111101000;
assign supra2[35][0] = 9'b111101000;
assign supra2[35][1] = 9'b111101000;
assign supra2[35][2] = 9'b111101000;
assign supra2[35][3] = 9'b101101000;
assign supra2[35][4] = 9'b100001111;
assign supra2[35][5] = 9'b100001111;
assign supra2[35][6] = 9'b100001111;
assign supra2[35][7] = 9'b100001111;
assign supra2[35][8] = 9'b100001111;
assign supra2[35][9] = 9'b100001111;
assign supra2[35][10] = 9'b100001111;
assign supra2[35][11] = 9'b100001111;
assign supra2[35][12] = 9'b100001111;
assign supra2[35][13] = 9'b100001111;
assign supra2[35][14] = 9'b101101000;
assign supra2[35][15] = 9'b111101000;
assign supra2[35][16] = 9'b111101000;
assign supra2[35][17] = 9'b111101000;
assign supra2[36][0] = 9'b111101000;
assign supra2[36][1] = 9'b111101000;
assign supra2[36][2] = 9'b111101000;
assign supra2[36][3] = 9'b101001001;
assign supra2[36][4] = 9'b100001111;
assign supra2[36][5] = 9'b100001111;
assign supra2[36][6] = 9'b100001111;
assign supra2[36][7] = 9'b100001111;
assign supra2[36][8] = 9'b100001111;
assign supra2[36][9] = 9'b100001111;
assign supra2[36][10] = 9'b100001111;
assign supra2[36][11] = 9'b100001111;
assign supra2[36][12] = 9'b100001111;
assign supra2[36][13] = 9'b100001111;
assign supra2[36][14] = 9'b101001001;
assign supra2[36][15] = 9'b111101000;
assign supra2[36][16] = 9'b111101000;
assign supra2[36][17] = 9'b111101000;
assign supra2[37][0] = 9'b111101000;
assign supra2[37][1] = 9'b111101000;
assign supra2[37][2] = 9'b111101000;
assign supra2[37][3] = 9'b101001000;
assign supra2[37][4] = 9'b100001111;
assign supra2[37][5] = 9'b100001111;
assign supra2[37][6] = 9'b100001111;
assign supra2[37][7] = 9'b100001111;
assign supra2[37][8] = 9'b100001111;
assign supra2[37][9] = 9'b100001111;
assign supra2[37][10] = 9'b100001111;
assign supra2[37][11] = 9'b100001111;
assign supra2[37][12] = 9'b100001111;
assign supra2[37][13] = 9'b100001111;
assign supra2[37][14] = 9'b101001001;
assign supra2[37][15] = 9'b111101000;
assign supra2[37][16] = 9'b111101000;
assign supra2[37][17] = 9'b111101000;
assign supra2[38][0] = 9'b111101000;
assign supra2[38][1] = 9'b111101000;
assign supra2[38][2] = 9'b111101000;
assign supra2[38][3] = 9'b110001000;
assign supra2[38][4] = 9'b100001010;
assign supra2[38][5] = 9'b100001111;
assign supra2[38][6] = 9'b100001111;
assign supra2[38][7] = 9'b100001111;
assign supra2[38][8] = 9'b100001111;
assign supra2[38][9] = 9'b100001111;
assign supra2[38][10] = 9'b100001111;
assign supra2[38][11] = 9'b100001111;
assign supra2[38][12] = 9'b100001111;
assign supra2[38][13] = 9'b100001010;
assign supra2[38][14] = 9'b110001000;
assign supra2[38][15] = 9'b111101000;
assign supra2[38][16] = 9'b111101000;
assign supra2[38][17] = 9'b111101000;
assign supra2[39][1] = 9'b111101000;
assign supra2[39][2] = 9'b111101000;
assign supra2[39][3] = 9'b111101000;
assign supra2[39][4] = 9'b110001000;
assign supra2[39][5] = 9'b100101001;
assign supra2[39][6] = 9'b100001010;
assign supra2[39][7] = 9'b100001111;
assign supra2[39][8] = 9'b100001111;
assign supra2[39][9] = 9'b100001111;
assign supra2[39][10] = 9'b100001111;
assign supra2[39][11] = 9'b100001010;
assign supra2[39][12] = 9'b100101001;
assign supra2[39][13] = 9'b110001000;
assign supra2[39][14] = 9'b111101000;
assign supra2[39][15] = 9'b111101000;
assign supra2[39][16] = 9'b111101000;
assign supra2[40][1] = 9'b111101000;
assign supra2[40][2] = 9'b111101000;
assign supra2[40][3] = 9'b111101000;
assign supra2[40][4] = 9'b111101000;
assign supra2[40][5] = 9'b111101000;
assign supra2[40][6] = 9'b111101000;
assign supra2[40][7] = 9'b110001000;
assign supra2[40][8] = 9'b110001000;
assign supra2[40][9] = 9'b110001000;
assign supra2[40][10] = 9'b110001000;
assign supra2[40][11] = 9'b111101000;
assign supra2[40][12] = 9'b111101000;
assign supra2[40][13] = 9'b111101000;
assign supra2[40][14] = 9'b111101000;
assign supra2[40][15] = 9'b111101000;
assign supra2[40][16] = 9'b111101000;
assign supra2[41][1] = 9'b111101000;
assign supra2[41][2] = 9'b111101000;
assign supra2[41][3] = 9'b110101000;
assign supra2[41][4] = 9'b110101000;
assign supra2[41][5] = 9'b111101000;
assign supra2[41][6] = 9'b111101000;
assign supra2[41][7] = 9'b111101000;
assign supra2[41][8] = 9'b111101000;
assign supra2[41][9] = 9'b111101000;
assign supra2[41][10] = 9'b111101000;
assign supra2[41][11] = 9'b111101000;
assign supra2[41][12] = 9'b111101000;
assign supra2[41][13] = 9'b110101000;
assign supra2[41][14] = 9'b110101000;
assign supra2[41][15] = 9'b111101000;
assign supra2[41][16] = 9'b111101000;
assign supra2[42][2] = 9'b110001000;
assign supra2[42][3] = 9'b101001101;
assign supra2[42][4] = 9'b101001101;
assign supra2[42][5] = 9'b101001101;
assign supra2[42][6] = 9'b101001101;
assign supra2[42][7] = 9'b101001101;
assign supra2[42][8] = 9'b101001101;
assign supra2[42][9] = 9'b101001101;
assign supra2[42][10] = 9'b101001101;
assign supra2[42][11] = 9'b101001101;
assign supra2[42][12] = 9'b101001101;
assign supra2[42][13] = 9'b101001101;
assign supra2[42][14] = 9'b101001101;
assign supra2[42][15] = 9'b110001000;
assign supra2[43][2] = 9'b101101000;
assign supra2[43][3] = 9'b101101101;
assign supra2[43][4] = 9'b101101101;
assign supra2[43][5] = 9'b101101101;
assign supra2[43][6] = 9'b101101101;
assign supra2[43][7] = 9'b101101101;
assign supra2[43][8] = 9'b101101101;
assign supra2[43][9] = 9'b101101101;
assign supra2[43][10] = 9'b101101101;
assign supra2[43][11] = 9'b101101101;
assign supra2[43][12] = 9'b101101101;
assign supra2[43][13] = 9'b101101101;
assign supra2[43][14] = 9'b101101101;
assign supra2[43][15] = 9'b101101000;
assign supra2[44][3] = 9'b111101000;
assign supra2[44][4] = 9'b111101000;
assign supra2[44][5] = 9'b111101000;
assign supra2[44][6] = 9'b111101000;
assign supra2[44][7] = 9'b111101000;
assign supra2[44][8] = 9'b111101000;
assign supra2[44][9] = 9'b111101000;
assign supra2[44][10] = 9'b111101000;
assign supra2[44][11] = 9'b111101000;
assign supra2[44][12] = 9'b111101000;
assign supra2[44][13] = 9'b111101000;
assign supra2[44][14] = 9'b110101000;
//Total de Lineas = 733
endmodule

