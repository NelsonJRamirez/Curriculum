`timescale 1ns / 1ps
module logo_rueda (
input enable,
input clock,
input [9:0] posx, posy,
input [9:0] hcount,
input [9:0] vcount,
output reg[2:0] red,
output reg[2:0] green,
output reg[1:0] blue,
output reg data);

always @(posedge clock)
begin
	if(enable)
	begin
		if(hcount >= posx & hcount < posx + RESOLUCION_X & vcount >= posy & vcount < posy + RESOLUCION_Y)
		begin
			if (logo_rueda[vcount - posy][hcount - posx][8] == 1'b1)
			begin
				red   <= logo_rueda[vcount- posy][hcount- posx][7:5];
				green <= logo_rueda[vcount- posy][hcount- posx][4:2];
            blue 	<= logo_rueda[vcount- posy][hcount- posx][1:0];
				data  <= 1'b1;
			end
			else
				data <= 0;
			end
		else
		data <= 0;
	end
end

parameter RESOLUCION_X = 50;
parameter RESOLUCION_Y = 50;
wire [8:0] logo_rueda[RESOLUCION_Y - 1'b1 : 0][RESOLUCION_X - 1'b1 : 0];
assign logo_rueda[1][8] = 9'b111101100;
assign logo_rueda[1][9] = 9'b111101100;
assign logo_rueda[1][10] = 9'b111100100;
assign logo_rueda[1][15] = 9'b110000100;
assign logo_rueda[1][16] = 9'b110101000;
assign logo_rueda[1][17] = 9'b111101000;
assign logo_rueda[1][18] = 9'b111101100;
assign logo_rueda[1][47] = 9'b101100100;
assign logo_rueda[1][48] = 9'b111101000;
assign logo_rueda[2][6] = 9'b111101100;
assign logo_rueda[2][7] = 9'b111101100;
assign logo_rueda[2][8] = 9'b111101100;
assign logo_rueda[2][9] = 9'b111101000;
assign logo_rueda[2][10] = 9'b111101000;
assign logo_rueda[2][11] = 9'b111101100;
assign logo_rueda[2][12] = 9'b111101100;
assign logo_rueda[2][13] = 9'b111101100;
assign logo_rueda[2][14] = 9'b111101100;
assign logo_rueda[2][15] = 9'b111101000;
assign logo_rueda[2][17] = 9'b101100100;
assign logo_rueda[2][18] = 9'b110000100;
assign logo_rueda[2][19] = 9'b111101000;
assign logo_rueda[2][20] = 9'b111101100;
assign logo_rueda[2][21] = 9'b111110000;
assign logo_rueda[2][47] = 9'b101000000;
assign logo_rueda[2][48] = 9'b110101000;
assign logo_rueda[3][4] = 9'b111101000;
assign logo_rueda[3][5] = 9'b111110000;
assign logo_rueda[3][6] = 9'b111110000;
assign logo_rueda[3][7] = 9'b111101000;
assign logo_rueda[3][8] = 9'b111101000;
assign logo_rueda[3][9] = 9'b111110000;
assign logo_rueda[3][10] = 9'b111111100;
assign logo_rueda[3][11] = 9'b111110100;
assign logo_rueda[3][12] = 9'b111101000;
assign logo_rueda[3][13] = 9'b111100100;
assign logo_rueda[3][19] = 9'b101000000;
assign logo_rueda[3][20] = 9'b110000100;
assign logo_rueda[3][21] = 9'b111110000;
assign logo_rueda[3][22] = 9'b111110000;
assign logo_rueda[3][23] = 9'b111110000;
assign logo_rueda[3][24] = 9'b111101100;
assign logo_rueda[3][46] = 9'b111101100;
assign logo_rueda[3][48] = 9'b111101100;
assign logo_rueda[4][3] = 9'b111101000;
assign logo_rueda[4][4] = 9'b111110000;
assign logo_rueda[4][5] = 9'b111110000;
assign logo_rueda[4][6] = 9'b111110000;
assign logo_rueda[4][7] = 9'b111110000;
assign logo_rueda[4][8] = 9'b111111100;
assign logo_rueda[4][9] = 9'b111111100;
assign logo_rueda[4][10] = 9'b111110100;
assign logo_rueda[4][11] = 9'b111110000;
assign logo_rueda[4][12] = 9'b111101100;
assign logo_rueda[4][13] = 9'b111110000;
assign logo_rueda[4][14] = 9'b111110000;
assign logo_rueda[4][15] = 9'b111110000;
assign logo_rueda[4][16] = 9'b111110000;
assign logo_rueda[4][17] = 9'b111110000;
assign logo_rueda[4][18] = 9'b111110000;
assign logo_rueda[4][19] = 9'b111110000;
assign logo_rueda[4][20] = 9'b110001000;
assign logo_rueda[4][21] = 9'b110000100;
assign logo_rueda[4][22] = 9'b111110000;
assign logo_rueda[4][23] = 9'b111110000;
assign logo_rueda[4][24] = 9'b111110000;
assign logo_rueda[4][25] = 9'b111110000;
assign logo_rueda[4][26] = 9'b111101100;
assign logo_rueda[4][45] = 9'b110101000;
assign logo_rueda[4][46] = 9'b111101100;
assign logo_rueda[4][47] = 9'b101100000;
assign logo_rueda[4][48] = 9'b111110000;
assign logo_rueda[5][3] = 9'b111110000;
assign logo_rueda[5][4] = 9'b111101000;
assign logo_rueda[5][5] = 9'b111101000;
assign logo_rueda[5][6] = 9'b111101100;
assign logo_rueda[5][7] = 9'b111111100;
assign logo_rueda[5][8] = 9'b111111100;
assign logo_rueda[5][9] = 9'b111110000;
assign logo_rueda[5][10] = 9'b111110000;
assign logo_rueda[5][11] = 9'b111110000;
assign logo_rueda[5][12] = 9'b111101000;
assign logo_rueda[5][13] = 9'b111101000;
assign logo_rueda[5][14] = 9'b111101000;
assign logo_rueda[5][15] = 9'b111101000;
assign logo_rueda[5][16] = 9'b111110000;
assign logo_rueda[5][17] = 9'b111101100;
assign logo_rueda[5][18] = 9'b111110000;
assign logo_rueda[5][19] = 9'b111101100;
assign logo_rueda[5][20] = 9'b111101100;
assign logo_rueda[5][21] = 9'b111110000;
assign logo_rueda[5][22] = 9'b111110100;
assign logo_rueda[5][23] = 9'b111101100;
assign logo_rueda[5][24] = 9'b111100100;
assign logo_rueda[5][25] = 9'b111101000;
assign logo_rueda[5][26] = 9'b111101100;
assign logo_rueda[5][27] = 9'b111110000;
assign logo_rueda[5][28] = 9'b111110000;
assign logo_rueda[5][29] = 9'b111101100;
assign logo_rueda[5][44] = 9'b110100100;
assign logo_rueda[5][45] = 9'b111110000;
assign logo_rueda[5][46] = 9'b111110000;
assign logo_rueda[5][47] = 9'b111110000;
assign logo_rueda[5][48] = 9'b111110100;
assign logo_rueda[6][2] = 9'b111101100;
assign logo_rueda[6][3] = 9'b111101100;
assign logo_rueda[6][4] = 9'b111100100;
assign logo_rueda[6][5] = 9'b111101000;
assign logo_rueda[6][6] = 9'b111101100;
assign logo_rueda[6][7] = 9'b111111100;
assign logo_rueda[6][8] = 9'b111111100;
assign logo_rueda[6][9] = 9'b111110000;
assign logo_rueda[6][10] = 9'b111110000;
assign logo_rueda[6][11] = 9'b111101000;
assign logo_rueda[6][12] = 9'b111100100;
assign logo_rueda[6][13] = 9'b111100100;
assign logo_rueda[6][14] = 9'b111101000;
assign logo_rueda[6][15] = 9'b111101100;
assign logo_rueda[6][16] = 9'b111110000;
assign logo_rueda[6][17] = 9'b111101100;
assign logo_rueda[6][18] = 9'b111101100;
assign logo_rueda[6][19] = 9'b111100100;
assign logo_rueda[6][20] = 9'b111100100;
assign logo_rueda[6][21] = 9'b111101000;
assign logo_rueda[6][22] = 9'b111101100;
assign logo_rueda[6][23] = 9'b111101100;
assign logo_rueda[6][24] = 9'b111101000;
assign logo_rueda[6][25] = 9'b111100100;
assign logo_rueda[6][26] = 9'b111100100;
assign logo_rueda[6][27] = 9'b111101000;
assign logo_rueda[6][28] = 9'b111101100;
assign logo_rueda[6][29] = 9'b111110000;
assign logo_rueda[6][30] = 9'b111110000;
assign logo_rueda[6][31] = 9'b111101100;
assign logo_rueda[6][43] = 9'b111101000;
assign logo_rueda[6][44] = 9'b111110000;
assign logo_rueda[6][45] = 9'b111110000;
assign logo_rueda[6][46] = 9'b111101000;
assign logo_rueda[6][47] = 9'b111101000;
assign logo_rueda[6][48] = 9'b111110000;
assign logo_rueda[7][1] = 9'b110000100;
assign logo_rueda[7][2] = 9'b111110000;
assign logo_rueda[7][3] = 9'b111101000;
assign logo_rueda[7][4] = 9'b111101000;
assign logo_rueda[7][5] = 9'b111101000;
assign logo_rueda[7][6] = 9'b111110000;
assign logo_rueda[7][7] = 9'b111111100;
assign logo_rueda[7][8] = 9'b111110000;
assign logo_rueda[7][9] = 9'b111110000;
assign logo_rueda[7][10] = 9'b111101100;
assign logo_rueda[7][11] = 9'b111101100;
assign logo_rueda[7][12] = 9'b111101100;
assign logo_rueda[7][13] = 9'b111101100;
assign logo_rueda[7][14] = 9'b111110000;
assign logo_rueda[7][15] = 9'b111110100;
assign logo_rueda[7][16] = 9'b111110000;
assign logo_rueda[7][17] = 9'b111110000;
assign logo_rueda[7][18] = 9'b111101000;
assign logo_rueda[7][19] = 9'b111100100;
assign logo_rueda[7][20] = 9'b111101000;
assign logo_rueda[7][21] = 9'b111101000;
assign logo_rueda[7][22] = 9'b111101000;
assign logo_rueda[7][23] = 9'b111101100;
assign logo_rueda[7][24] = 9'b111101000;
assign logo_rueda[7][25] = 9'b111101000;
assign logo_rueda[7][26] = 9'b111100100;
assign logo_rueda[7][27] = 9'b111101000;
assign logo_rueda[7][28] = 9'b111101000;
assign logo_rueda[7][29] = 9'b111101000;
assign logo_rueda[7][30] = 9'b111101100;
assign logo_rueda[7][31] = 9'b111110000;
assign logo_rueda[7][32] = 9'b111110000;
assign logo_rueda[7][33] = 9'b111110000;
assign logo_rueda[7][34] = 9'b111110000;
assign logo_rueda[7][35] = 9'b111101100;
assign logo_rueda[7][36] = 9'b111101100;
assign logo_rueda[7][41] = 9'b111101100;
assign logo_rueda[7][42] = 9'b111110000;
assign logo_rueda[7][43] = 9'b111110100;
assign logo_rueda[7][44] = 9'b111110000;
assign logo_rueda[7][45] = 9'b111110000;
assign logo_rueda[7][46] = 9'b111101000;
assign logo_rueda[7][47] = 9'b111100100;
assign logo_rueda[7][48] = 9'b111110000;
assign logo_rueda[8][1] = 9'b110101000;
assign logo_rueda[8][2] = 9'b111101100;
assign logo_rueda[8][3] = 9'b111101000;
assign logo_rueda[8][4] = 9'b111101000;
assign logo_rueda[8][5] = 9'b111101000;
assign logo_rueda[8][6] = 9'b111101100;
assign logo_rueda[8][7] = 9'b111110000;
assign logo_rueda[8][8] = 9'b111110000;
assign logo_rueda[8][9] = 9'b111101100;
assign logo_rueda[8][10] = 9'b111110000;
assign logo_rueda[8][11] = 9'b111110100;
assign logo_rueda[8][12] = 9'b111110000;
assign logo_rueda[8][13] = 9'b111101100;
assign logo_rueda[8][14] = 9'b111101100;
assign logo_rueda[8][15] = 9'b111110000;
assign logo_rueda[8][16] = 9'b111110000;
assign logo_rueda[8][17] = 9'b111110100;
assign logo_rueda[8][18] = 9'b111101100;
assign logo_rueda[8][19] = 9'b111101000;
assign logo_rueda[8][20] = 9'b111101000;
assign logo_rueda[8][21] = 9'b111101000;
assign logo_rueda[8][22] = 9'b111101000;
assign logo_rueda[8][23] = 9'b111101100;
assign logo_rueda[8][24] = 9'b111101100;
assign logo_rueda[8][25] = 9'b111101100;
assign logo_rueda[8][26] = 9'b111101000;
assign logo_rueda[8][27] = 9'b111101000;
assign logo_rueda[8][28] = 9'b111101000;
assign logo_rueda[8][29] = 9'b111101000;
assign logo_rueda[8][30] = 9'b111101000;
assign logo_rueda[8][31] = 9'b111101000;
assign logo_rueda[8][32] = 9'b111101000;
assign logo_rueda[8][33] = 9'b111101100;
assign logo_rueda[8][34] = 9'b111110000;
assign logo_rueda[8][35] = 9'b111110000;
assign logo_rueda[8][36] = 9'b111110000;
assign logo_rueda[8][37] = 9'b111110000;
assign logo_rueda[8][38] = 9'b111110000;
assign logo_rueda[8][39] = 9'b111110000;
assign logo_rueda[8][40] = 9'b111110100;
assign logo_rueda[8][41] = 9'b111110100;
assign logo_rueda[8][42] = 9'b111110000;
assign logo_rueda[8][43] = 9'b111101100;
assign logo_rueda[8][44] = 9'b111101100;
assign logo_rueda[8][45] = 9'b111110000;
assign logo_rueda[8][46] = 9'b111110100;
assign logo_rueda[8][47] = 9'b111110000;
assign logo_rueda[8][48] = 9'b111110000;
assign logo_rueda[9][1] = 9'b111101100;
assign logo_rueda[9][2] = 9'b111101100;
assign logo_rueda[9][3] = 9'b111101000;
assign logo_rueda[9][4] = 9'b111101000;
assign logo_rueda[9][5] = 9'b111101000;
assign logo_rueda[9][6] = 9'b111101000;
assign logo_rueda[9][7] = 9'b111110000;
assign logo_rueda[9][8] = 9'b111110000;
assign logo_rueda[9][9] = 9'b111110100;
assign logo_rueda[9][10] = 9'b111110100;
assign logo_rueda[9][11] = 9'b110001100;
assign logo_rueda[9][12] = 9'b101101000;
assign logo_rueda[9][13] = 9'b101000100;
assign logo_rueda[9][14] = 9'b100100100;
assign logo_rueda[9][15] = 9'b101000100;
assign logo_rueda[9][16] = 9'b101000100;
assign logo_rueda[9][17] = 9'b110001000;
assign logo_rueda[9][18] = 9'b111101100;
assign logo_rueda[9][19] = 9'b111110000;
assign logo_rueda[9][20] = 9'b111101100;
assign logo_rueda[9][21] = 9'b111101000;
assign logo_rueda[9][22] = 9'b111101000;
assign logo_rueda[9][23] = 9'b111101100;
assign logo_rueda[9][24] = 9'b111101100;
assign logo_rueda[9][25] = 9'b111101100;
assign logo_rueda[9][26] = 9'b111101000;
assign logo_rueda[9][27] = 9'b111101000;
assign logo_rueda[9][28] = 9'b111101000;
assign logo_rueda[9][29] = 9'b111101000;
assign logo_rueda[9][30] = 9'b111101000;
assign logo_rueda[9][31] = 9'b111101000;
assign logo_rueda[9][32] = 9'b111101000;
assign logo_rueda[9][33] = 9'b111101000;
assign logo_rueda[9][34] = 9'b111101000;
assign logo_rueda[9][35] = 9'b111101000;
assign logo_rueda[9][36] = 9'b111101100;
assign logo_rueda[9][37] = 9'b111101100;
assign logo_rueda[9][38] = 9'b111110000;
assign logo_rueda[9][39] = 9'b111110000;
assign logo_rueda[9][40] = 9'b111110000;
assign logo_rueda[9][41] = 9'b111110000;
assign logo_rueda[9][42] = 9'b111101100;
assign logo_rueda[9][43] = 9'b111101100;
assign logo_rueda[9][44] = 9'b111101100;
assign logo_rueda[9][45] = 9'b111110000;
assign logo_rueda[9][46] = 9'b111110100;
assign logo_rueda[9][47] = 9'b111101000;
assign logo_rueda[9][48] = 9'b111110000;
assign logo_rueda[10][1] = 9'b111101100;
assign logo_rueda[10][2] = 9'b111101100;
assign logo_rueda[10][3] = 9'b111101100;
assign logo_rueda[10][4] = 9'b111101100;
assign logo_rueda[10][5] = 9'b111101000;
assign logo_rueda[10][6] = 9'b111110000;
assign logo_rueda[10][7] = 9'b111110100;
assign logo_rueda[10][8] = 9'b111110100;
assign logo_rueda[10][9] = 9'b111110100;
assign logo_rueda[10][10] = 9'b101101000;
assign logo_rueda[10][11] = 9'b100101001;
assign logo_rueda[10][12] = 9'b100100100;
assign logo_rueda[10][13] = 9'b101001000;
assign logo_rueda[10][14] = 9'b101101100;
assign logo_rueda[10][15] = 9'b101101100;
assign logo_rueda[10][16] = 9'b100101000;
assign logo_rueda[10][17] = 9'b100100100;
assign logo_rueda[10][18] = 9'b100100100;
assign logo_rueda[10][19] = 9'b101100100;
assign logo_rueda[10][20] = 9'b111101100;
assign logo_rueda[10][21] = 9'b111110000;
assign logo_rueda[10][22] = 9'b111101100;
assign logo_rueda[10][23] = 9'b111101100;
assign logo_rueda[10][24] = 9'b111101100;
assign logo_rueda[10][25] = 9'b111101100;
assign logo_rueda[10][26] = 9'b111101100;
assign logo_rueda[10][27] = 9'b111101000;
assign logo_rueda[10][28] = 9'b111101000;
assign logo_rueda[10][29] = 9'b111101000;
assign logo_rueda[10][30] = 9'b111101000;
assign logo_rueda[10][31] = 9'b111101000;
assign logo_rueda[10][32] = 9'b111101000;
assign logo_rueda[10][33] = 9'b111101000;
assign logo_rueda[10][34] = 9'b111101000;
assign logo_rueda[10][35] = 9'b111101100;
assign logo_rueda[10][36] = 9'b111101100;
assign logo_rueda[10][37] = 9'b111101100;
assign logo_rueda[10][38] = 9'b111101100;
assign logo_rueda[10][39] = 9'b111101100;
assign logo_rueda[10][40] = 9'b111101100;
assign logo_rueda[10][41] = 9'b111110000;
assign logo_rueda[10][42] = 9'b111110000;
assign logo_rueda[10][43] = 9'b111110000;
assign logo_rueda[10][44] = 9'b111110100;
assign logo_rueda[10][45] = 9'b111110100;
assign logo_rueda[10][46] = 9'b111110000;
assign logo_rueda[10][47] = 9'b110000100;
assign logo_rueda[10][48] = 9'b111110000;
assign logo_rueda[11][1] = 9'b111101100;
assign logo_rueda[11][2] = 9'b111110000;
assign logo_rueda[11][3] = 9'b111110000;
assign logo_rueda[11][4] = 9'b111101100;
assign logo_rueda[11][5] = 9'b111101100;
assign logo_rueda[11][6] = 9'b111110000;
assign logo_rueda[11][7] = 9'b111101100;
assign logo_rueda[11][8] = 9'b111111100;
assign logo_rueda[11][9] = 9'b110001000;
assign logo_rueda[11][10] = 9'b100101001;
assign logo_rueda[11][11] = 9'b100100100;
assign logo_rueda[11][12] = 9'b111101100;
assign logo_rueda[11][13] = 9'b111111100;
assign logo_rueda[11][14] = 9'b111111100;
assign logo_rueda[11][15] = 9'b111111100;
assign logo_rueda[11][16] = 9'b111111101;
assign logo_rueda[11][17] = 9'b110010001;
assign logo_rueda[11][18] = 9'b101001000;
assign logo_rueda[11][19] = 9'b100100100;
assign logo_rueda[11][20] = 9'b101000100;
assign logo_rueda[11][21] = 9'b110001000;
assign logo_rueda[11][22] = 9'b111110000;
assign logo_rueda[11][23] = 9'b111110000;
assign logo_rueda[11][24] = 9'b111101100;
assign logo_rueda[11][25] = 9'b111101100;
assign logo_rueda[11][26] = 9'b111101100;
assign logo_rueda[11][27] = 9'b111101100;
assign logo_rueda[11][28] = 9'b111101100;
assign logo_rueda[11][29] = 9'b111101100;
assign logo_rueda[11][30] = 9'b111101100;
assign logo_rueda[11][31] = 9'b111101100;
assign logo_rueda[11][32] = 9'b111101100;
assign logo_rueda[11][33] = 9'b111101000;
assign logo_rueda[11][34] = 9'b111101100;
assign logo_rueda[11][35] = 9'b111101100;
assign logo_rueda[11][36] = 9'b111101100;
assign logo_rueda[11][37] = 9'b111101100;
assign logo_rueda[11][38] = 9'b111110000;
assign logo_rueda[11][39] = 9'b111101100;
assign logo_rueda[11][40] = 9'b111101100;
assign logo_rueda[11][41] = 9'b111110000;
assign logo_rueda[11][42] = 9'b111111100;
assign logo_rueda[11][43] = 9'b111110000;
assign logo_rueda[11][44] = 9'b111110000;
assign logo_rueda[11][45] = 9'b111111100;
assign logo_rueda[11][46] = 9'b111110000;
assign logo_rueda[11][47] = 9'b110000100;
assign logo_rueda[11][48] = 9'b111101100;
assign logo_rueda[12][0] = 9'b101000000;
assign logo_rueda[12][1] = 9'b111110000;
assign logo_rueda[12][2] = 9'b111110100;
assign logo_rueda[12][3] = 9'b111110000;
assign logo_rueda[12][4] = 9'b111110000;
assign logo_rueda[12][5] = 9'b111110000;
assign logo_rueda[12][6] = 9'b110101000;
assign logo_rueda[12][7] = 9'b111101100;
assign logo_rueda[12][8] = 9'b111110000;
assign logo_rueda[12][9] = 9'b101001001;
assign logo_rueda[12][10] = 9'b100101001;
assign logo_rueda[12][11] = 9'b101101000;
assign logo_rueda[12][12] = 9'b111110000;
assign logo_rueda[12][13] = 9'b111110000;
assign logo_rueda[12][14] = 9'b110101100;
assign logo_rueda[12][15] = 9'b110001000;
assign logo_rueda[12][16] = 9'b101101000;
assign logo_rueda[12][17] = 9'b110110000;
assign logo_rueda[12][18] = 9'b111111101;
assign logo_rueda[12][19] = 9'b110110001;
assign logo_rueda[12][20] = 9'b101001001;
assign logo_rueda[12][21] = 9'b100100100;
assign logo_rueda[12][22] = 9'b101100100;
assign logo_rueda[12][23] = 9'b111110000;
assign logo_rueda[12][24] = 9'b111110000;
assign logo_rueda[12][25] = 9'b111101100;
assign logo_rueda[12][26] = 9'b111101100;
assign logo_rueda[12][27] = 9'b111101100;
assign logo_rueda[12][28] = 9'b111101100;
assign logo_rueda[12][29] = 9'b111101100;
assign logo_rueda[12][30] = 9'b111101100;
assign logo_rueda[12][31] = 9'b111101100;
assign logo_rueda[12][32] = 9'b111101100;
assign logo_rueda[12][33] = 9'b111101100;
assign logo_rueda[12][34] = 9'b111101100;
assign logo_rueda[12][35] = 9'b111101100;
assign logo_rueda[12][36] = 9'b111110000;
assign logo_rueda[12][37] = 9'b111110000;
assign logo_rueda[12][38] = 9'b111110100;
assign logo_rueda[12][39] = 9'b111110100;
assign logo_rueda[12][40] = 9'b111110100;
assign logo_rueda[12][41] = 9'b111111100;
assign logo_rueda[12][42] = 9'b111110000;
assign logo_rueda[12][43] = 9'b101100000;
assign logo_rueda[12][44] = 9'b111110000;
assign logo_rueda[12][45] = 9'b111111100;
assign logo_rueda[12][47] = 9'b110101000;
assign logo_rueda[12][48] = 9'b111101100;
assign logo_rueda[13][1] = 9'b111110000;
assign logo_rueda[13][2] = 9'b111110000;
assign logo_rueda[13][3] = 9'b110001000;
assign logo_rueda[13][4] = 9'b111110000;
assign logo_rueda[13][5] = 9'b111110000;
assign logo_rueda[13][6] = 9'b110000100;
assign logo_rueda[13][7] = 9'b111110000;
assign logo_rueda[13][8] = 9'b111110000;
assign logo_rueda[13][9] = 9'b101001001;
assign logo_rueda[13][10] = 9'b101001001;
assign logo_rueda[13][11] = 9'b110101000;
assign logo_rueda[13][12] = 9'b111101100;
assign logo_rueda[13][13] = 9'b111101100;
assign logo_rueda[13][14] = 9'b110101001;
assign logo_rueda[13][15] = 9'b110001001;
assign logo_rueda[13][16] = 9'b101100100;
assign logo_rueda[13][17] = 9'b101000000;
assign logo_rueda[13][18] = 9'b101100100;
assign logo_rueda[13][19] = 9'b110001100;
assign logo_rueda[13][20] = 9'b111110001;
assign logo_rueda[13][21] = 9'b101101101;
assign logo_rueda[13][22] = 9'b100100100;
assign logo_rueda[13][23] = 9'b101100100;
assign logo_rueda[13][24] = 9'b111110000;
assign logo_rueda[13][25] = 9'b111110100;
assign logo_rueda[13][26] = 9'b111110100;
assign logo_rueda[13][27] = 9'b111101100;
assign logo_rueda[13][28] = 9'b111101100;
assign logo_rueda[13][29] = 9'b111101100;
assign logo_rueda[13][30] = 9'b111101100;
assign logo_rueda[13][31] = 9'b111110100;
assign logo_rueda[13][32] = 9'b111110000;
assign logo_rueda[13][33] = 9'b111110000;
assign logo_rueda[13][34] = 9'b111110000;
assign logo_rueda[13][35] = 9'b111110000;
assign logo_rueda[13][36] = 9'b111111100;
assign logo_rueda[13][37] = 9'b111110000;
assign logo_rueda[13][38] = 9'b111101100;
assign logo_rueda[13][39] = 9'b111101100;
assign logo_rueda[13][40] = 9'b111101100;
assign logo_rueda[13][41] = 9'b111101000;
assign logo_rueda[13][44] = 9'b111110100;
assign logo_rueda[13][45] = 9'b111110000;
assign logo_rueda[13][46] = 9'b110100100;
assign logo_rueda[13][47] = 9'b111101000;
assign logo_rueda[14][1] = 9'b111101100;
assign logo_rueda[14][2] = 9'b111110000;
assign logo_rueda[14][3] = 9'b110001000;
assign logo_rueda[14][4] = 9'b111110100;
assign logo_rueda[14][5] = 9'b111110000;
assign logo_rueda[14][6] = 9'b101100000;
assign logo_rueda[14][7] = 9'b111110000;
assign logo_rueda[14][8] = 9'b110101100;
assign logo_rueda[14][9] = 9'b101001001;
assign logo_rueda[14][10] = 9'b101001001;
assign logo_rueda[14][11] = 9'b110101100;
assign logo_rueda[14][12] = 9'b111101000;
assign logo_rueda[14][13] = 9'b111101101;
assign logo_rueda[14][14] = 9'b111111111;
assign logo_rueda[14][15] = 9'b111111111;
assign logo_rueda[14][16] = 9'b111110001;
assign logo_rueda[14][17] = 9'b111101101;
assign logo_rueda[14][18] = 9'b110101001;
assign logo_rueda[14][19] = 9'b110000100;
assign logo_rueda[14][20] = 9'b101100100;
assign logo_rueda[14][21] = 9'b111101100;
assign logo_rueda[14][22] = 9'b110001101;
assign logo_rueda[14][23] = 9'b100100101;
assign logo_rueda[14][24] = 9'b101100100;
assign logo_rueda[14][25] = 9'b111110000;
assign logo_rueda[14][26] = 9'b111110000;
assign logo_rueda[14][27] = 9'b111110000;
assign logo_rueda[14][28] = 9'b111110000;
assign logo_rueda[14][29] = 9'b111110000;
assign logo_rueda[14][30] = 9'b111110000;
assign logo_rueda[14][31] = 9'b111110100;
assign logo_rueda[14][32] = 9'b110101100;
assign logo_rueda[14][33] = 9'b110000100;
assign logo_rueda[14][34] = 9'b110101100;
assign logo_rueda[14][35] = 9'b111110000;
assign logo_rueda[14][36] = 9'b111110100;
assign logo_rueda[14][37] = 9'b111110000;
assign logo_rueda[14][38] = 9'b111101100;
assign logo_rueda[14][39] = 9'b111101000;
assign logo_rueda[14][40] = 9'b111101000;
assign logo_rueda[14][43] = 9'b111101100;
assign logo_rueda[14][44] = 9'b111101100;
assign logo_rueda[15][1] = 9'b110101000;
assign logo_rueda[15][2] = 9'b111110000;
assign logo_rueda[15][3] = 9'b110000100;
assign logo_rueda[15][4] = 9'b111111100;
assign logo_rueda[15][5] = 9'b111110000;
assign logo_rueda[15][6] = 9'b101100000;
assign logo_rueda[15][7] = 9'b111110000;
assign logo_rueda[15][8] = 9'b110101100;
assign logo_rueda[15][9] = 9'b101001001;
assign logo_rueda[15][10] = 9'b100101001;
assign logo_rueda[15][11] = 9'b110001000;
assign logo_rueda[15][12] = 9'b111101000;
assign logo_rueda[15][13] = 9'b111101101;
assign logo_rueda[15][14] = 9'b111111111;
assign logo_rueda[15][15] = 9'b111111111;
assign logo_rueda[15][16] = 9'b111111111;
assign logo_rueda[15][17] = 9'b111111111;
assign logo_rueda[15][18] = 9'b111110101;
assign logo_rueda[15][19] = 9'b111110001;
assign logo_rueda[15][20] = 9'b111101000;
assign logo_rueda[15][21] = 9'b110000100;
assign logo_rueda[15][22] = 9'b111101100;
assign logo_rueda[15][23] = 9'b110001101;
assign logo_rueda[15][24] = 9'b100101001;
assign logo_rueda[15][25] = 9'b101100100;
assign logo_rueda[15][26] = 9'b110101000;
assign logo_rueda[15][27] = 9'b110000100;
assign logo_rueda[15][28] = 9'b111110100;
assign logo_rueda[15][29] = 9'b111110100;
assign logo_rueda[15][30] = 9'b111110000;
assign logo_rueda[15][31] = 9'b111110000;
assign logo_rueda[15][32] = 9'b111110100;
assign logo_rueda[15][33] = 9'b111110000;
assign logo_rueda[15][34] = 9'b110000100;
assign logo_rueda[15][35] = 9'b110000100;
assign logo_rueda[15][36] = 9'b110000100;
assign logo_rueda[15][37] = 9'b110001000;
assign logo_rueda[15][38] = 9'b110101000;
assign logo_rueda[15][39] = 9'b111101100;
assign logo_rueda[15][40] = 9'b111101100;
assign logo_rueda[15][42] = 9'b111101000;
assign logo_rueda[15][43] = 9'b111101000;
assign logo_rueda[16][1] = 9'b110000100;
assign logo_rueda[16][2] = 9'b111110000;
assign logo_rueda[16][3] = 9'b101100000;
assign logo_rueda[16][4] = 9'b111110100;
assign logo_rueda[16][5] = 9'b111110100;
assign logo_rueda[16][6] = 9'b101000000;
assign logo_rueda[16][7] = 9'b111110000;
assign logo_rueda[16][8] = 9'b111110000;
assign logo_rueda[16][9] = 9'b101001001;
assign logo_rueda[16][10] = 9'b101001001;
assign logo_rueda[16][11] = 9'b101101000;
assign logo_rueda[16][12] = 9'b111101000;
assign logo_rueda[16][13] = 9'b111101101;
assign logo_rueda[16][14] = 9'b111110001;
assign logo_rueda[16][15] = 9'b111111110;
assign logo_rueda[16][16] = 9'b111111111;
assign logo_rueda[16][17] = 9'b111110001;
assign logo_rueda[16][18] = 9'b110100100;
assign logo_rueda[16][19] = 9'b111110000;
assign logo_rueda[16][20] = 9'b111110000;
assign logo_rueda[16][21] = 9'b110100100;
assign logo_rueda[16][22] = 9'b110000100;
assign logo_rueda[16][23] = 9'b111101000;
assign logo_rueda[16][24] = 9'b101101101;
assign logo_rueda[16][25] = 9'b100101001;
assign logo_rueda[16][26] = 9'b110001000;
assign logo_rueda[16][27] = 9'b101101000;
assign logo_rueda[16][28] = 9'b101100100;
assign logo_rueda[16][29] = 9'b111111100;
assign logo_rueda[16][30] = 9'b111111100;
assign logo_rueda[16][31] = 9'b111110100;
assign logo_rueda[16][32] = 9'b111110100;
assign logo_rueda[16][33] = 9'b111111100;
assign logo_rueda[16][34] = 9'b111111100;
assign logo_rueda[16][35] = 9'b111110000;
assign logo_rueda[16][42] = 9'b111100100;
assign logo_rueda[17][1] = 9'b101000000;
assign logo_rueda[17][2] = 9'b111101100;
assign logo_rueda[17][3] = 9'b101000000;
assign logo_rueda[17][4] = 9'b111110000;
assign logo_rueda[17][5] = 9'b111110100;
assign logo_rueda[17][6] = 9'b101000000;
assign logo_rueda[17][7] = 9'b110101100;
assign logo_rueda[17][8] = 9'b111110100;
assign logo_rueda[17][9] = 9'b101101001;
assign logo_rueda[17][10] = 9'b101001001;
assign logo_rueda[17][11] = 9'b101000100;
assign logo_rueda[17][12] = 9'b111101000;
assign logo_rueda[17][13] = 9'b111110001;
assign logo_rueda[17][14] = 9'b111110001;
assign logo_rueda[17][15] = 9'b111110001;
assign logo_rueda[17][16] = 9'b111111110;
assign logo_rueda[17][17] = 9'b111101001;
assign logo_rueda[17][18] = 9'b110001001;
assign logo_rueda[17][19] = 9'b111100100;
assign logo_rueda[17][20] = 9'b111101100;
assign logo_rueda[17][21] = 9'b111101000;
assign logo_rueda[17][22] = 9'b111110001;
assign logo_rueda[17][23] = 9'b111101101;
assign logo_rueda[17][24] = 9'b111101000;
assign logo_rueda[17][25] = 9'b101101101;
assign logo_rueda[17][26] = 9'b101001000;
assign logo_rueda[17][27] = 9'b110001000;
assign logo_rueda[17][28] = 9'b101000100;
assign logo_rueda[17][29] = 9'b110000100;
assign logo_rueda[17][30] = 9'b111110100;
assign logo_rueda[17][31] = 9'b111101100;
assign logo_rueda[17][32] = 9'b111110100;
assign logo_rueda[17][33] = 9'b111111100;
assign logo_rueda[17][34] = 9'b111111100;
assign logo_rueda[17][35] = 9'b111101100;
assign logo_rueda[17][37] = 9'b111101100;
assign logo_rueda[17][38] = 9'b111110000;
assign logo_rueda[17][39] = 9'b111110000;
assign logo_rueda[17][40] = 9'b111110000;
assign logo_rueda[17][41] = 9'b111110100;
assign logo_rueda[17][42] = 9'b111110000;
assign logo_rueda[17][43] = 9'b111101100;
assign logo_rueda[17][44] = 9'b111101000;
assign logo_rueda[18][2] = 9'b110001000;
assign logo_rueda[18][3] = 9'b101100100;
assign logo_rueda[18][4] = 9'b110101100;
assign logo_rueda[18][5] = 9'b111111100;
assign logo_rueda[18][6] = 9'b110000101;
assign logo_rueda[18][7] = 9'b110001000;
assign logo_rueda[18][8] = 9'b111111100;
assign logo_rueda[18][9] = 9'b101101001;
assign logo_rueda[18][10] = 9'b101001001;
assign logo_rueda[18][11] = 9'b100100100;
assign logo_rueda[18][12] = 9'b110101000;
assign logo_rueda[18][13] = 9'b111110001;
assign logo_rueda[18][14] = 9'b111111111;
assign logo_rueda[18][15] = 9'b111110101;
assign logo_rueda[18][16] = 9'b111110001;
assign logo_rueda[18][17] = 9'b111101000;
assign logo_rueda[18][18] = 9'b111110110;
assign logo_rueda[18][19] = 9'b111110001;
assign logo_rueda[18][20] = 9'b111100100;
assign logo_rueda[18][21] = 9'b111100100;
assign logo_rueda[18][22] = 9'b111111110;
assign logo_rueda[18][23] = 9'b111111111;
assign logo_rueda[18][24] = 9'b111100100;
assign logo_rueda[18][25] = 9'b111101000;
assign logo_rueda[18][26] = 9'b101001001;
assign logo_rueda[18][27] = 9'b101001001;
assign logo_rueda[18][28] = 9'b101101101;
assign logo_rueda[18][29] = 9'b100100100;
assign logo_rueda[18][30] = 9'b110000100;
assign logo_rueda[18][31] = 9'b111110000;
assign logo_rueda[18][32] = 9'b110101000;
assign logo_rueda[18][33] = 9'b111111100;
assign logo_rueda[18][34] = 9'b111111100;
assign logo_rueda[18][35] = 9'b111101100;
assign logo_rueda[18][36] = 9'b111110000;
assign logo_rueda[18][37] = 9'b111111100;
assign logo_rueda[18][38] = 9'b111111100;
assign logo_rueda[18][39] = 9'b111111100;
assign logo_rueda[18][40] = 9'b111111100;
assign logo_rueda[18][41] = 9'b111110100;
assign logo_rueda[18][42] = 9'b111101000;
assign logo_rueda[19][2] = 9'b101100100;
assign logo_rueda[19][3] = 9'b110001000;
assign logo_rueda[19][4] = 9'b110000100;
assign logo_rueda[19][5] = 9'b111111100;
assign logo_rueda[19][6] = 9'b111110001;
assign logo_rueda[19][7] = 9'b101000000;
assign logo_rueda[19][8] = 9'b111110100;
assign logo_rueda[19][9] = 9'b110001101;
assign logo_rueda[19][10] = 9'b101001001;
assign logo_rueda[19][11] = 9'b101001001;
assign logo_rueda[19][12] = 9'b101100100;
assign logo_rueda[19][13] = 9'b111101100;
assign logo_rueda[19][14] = 9'b111111111;
assign logo_rueda[19][15] = 9'b111111111;
assign logo_rueda[19][16] = 9'b111110001;
assign logo_rueda[19][17] = 9'b111101000;
assign logo_rueda[19][18] = 9'b110101101;
assign logo_rueda[19][19] = 9'b111111111;
assign logo_rueda[19][20] = 9'b111101101;
assign logo_rueda[19][21] = 9'b111100000;
assign logo_rueda[19][22] = 9'b111110001;
assign logo_rueda[19][23] = 9'b111111111;
assign logo_rueda[19][24] = 9'b111101000;
assign logo_rueda[19][25] = 9'b111101100;
assign logo_rueda[19][26] = 9'b110101101;
assign logo_rueda[19][27] = 9'b100100100;
assign logo_rueda[19][28] = 9'b101001001;
assign logo_rueda[19][29] = 9'b101001101;
assign logo_rueda[19][30] = 9'b100100100;
assign logo_rueda[19][31] = 9'b110001000;
assign logo_rueda[19][32] = 9'b111101100;
assign logo_rueda[19][33] = 9'b110101000;
assign logo_rueda[19][34] = 9'b111111100;
assign logo_rueda[19][35] = 9'b111111100;
assign logo_rueda[19][36] = 9'b111111100;
assign logo_rueda[19][37] = 9'b111111100;
assign logo_rueda[19][38] = 9'b111110100;
assign logo_rueda[19][39] = 9'b111111100;
assign logo_rueda[19][40] = 9'b111111100;
assign logo_rueda[19][41] = 9'b111110000;
assign logo_rueda[19][42] = 9'b111101100;
assign logo_rueda[19][43] = 9'b111101000;
assign logo_rueda[20][3] = 9'b110000100;
assign logo_rueda[20][4] = 9'b101000000;
assign logo_rueda[20][5] = 9'b111110100;
assign logo_rueda[20][6] = 9'b111110101;
assign logo_rueda[20][8] = 9'b111101100;
assign logo_rueda[20][9] = 9'b111110000;
assign logo_rueda[20][10] = 9'b101101001;
assign logo_rueda[20][11] = 9'b101001001;
assign logo_rueda[20][12] = 9'b100100100;
assign logo_rueda[20][13] = 9'b111101000;
assign logo_rueda[20][14] = 9'b111111110;
assign logo_rueda[20][15] = 9'b111111111;
assign logo_rueda[20][16] = 9'b111111110;
assign logo_rueda[20][17] = 9'b111101100;
assign logo_rueda[20][18] = 9'b111101000;
assign logo_rueda[20][19] = 9'b111101101;
assign logo_rueda[20][20] = 9'b111111110;
assign logo_rueda[20][21] = 9'b111101001;
assign logo_rueda[20][22] = 9'b111101101;
assign logo_rueda[20][23] = 9'b111110101;
assign logo_rueda[20][24] = 9'b111101000;
assign logo_rueda[20][25] = 9'b111111100;
assign logo_rueda[20][26] = 9'b111110100;
assign logo_rueda[20][27] = 9'b101101000;
assign logo_rueda[20][28] = 9'b100100100;
assign logo_rueda[20][29] = 9'b101101101;
assign logo_rueda[20][30] = 9'b101001001;
assign logo_rueda[20][31] = 9'b100100000;
assign logo_rueda[20][32] = 9'b111101100;
assign logo_rueda[20][33] = 9'b110001000;
assign logo_rueda[20][34] = 9'b111101100;
assign logo_rueda[20][35] = 9'b111111100;
assign logo_rueda[20][36] = 9'b111111100;
assign logo_rueda[20][37] = 9'b111111100;
assign logo_rueda[20][38] = 9'b111111100;
assign logo_rueda[20][39] = 9'b111111100;
assign logo_rueda[20][40] = 9'b111110000;
assign logo_rueda[20][41] = 9'b111101100;
assign logo_rueda[20][42] = 9'b111101000;
assign logo_rueda[20][43] = 9'b111101000;
assign logo_rueda[21][5] = 9'b110001000;
assign logo_rueda[21][6] = 9'b111110100;
assign logo_rueda[21][8] = 9'b101100100;
assign logo_rueda[21][9] = 9'b111111100;
assign logo_rueda[21][10] = 9'b110001101;
assign logo_rueda[21][11] = 9'b101001001;
assign logo_rueda[21][12] = 9'b101001001;
assign logo_rueda[21][13] = 9'b101100100;
assign logo_rueda[21][14] = 9'b111101100;
assign logo_rueda[21][15] = 9'b111111111;
assign logo_rueda[21][16] = 9'b111111110;
assign logo_rueda[21][17] = 9'b111110001;
assign logo_rueda[21][18] = 9'b111110000;
assign logo_rueda[21][19] = 9'b111101100;
assign logo_rueda[21][20] = 9'b111101101;
assign logo_rueda[21][21] = 9'b111110001;
assign logo_rueda[21][22] = 9'b111111111;
assign logo_rueda[21][23] = 9'b111110001;
assign logo_rueda[21][24] = 9'b111101000;
assign logo_rueda[21][25] = 9'b111111100;
assign logo_rueda[21][26] = 9'b111111100;
assign logo_rueda[21][27] = 9'b111110000;
assign logo_rueda[21][28] = 9'b100100100;
assign logo_rueda[21][29] = 9'b101001001;
assign logo_rueda[21][30] = 9'b101101101;
assign logo_rueda[21][31] = 9'b101001001;
assign logo_rueda[21][32] = 9'b101000000;
assign logo_rueda[21][33] = 9'b111101100;
assign logo_rueda[21][34] = 9'b101100100;
assign logo_rueda[21][35] = 9'b111110100;
assign logo_rueda[21][36] = 9'b111111100;
assign logo_rueda[21][37] = 9'b111111100;
assign logo_rueda[21][38] = 9'b111111100;
assign logo_rueda[21][39] = 9'b111110000;
assign logo_rueda[22][5] = 9'b101100000;
assign logo_rueda[22][6] = 9'b111110100;
assign logo_rueda[22][7] = 9'b111110001;
assign logo_rueda[22][8] = 9'b100100000;
assign logo_rueda[22][9] = 9'b111110000;
assign logo_rueda[22][10] = 9'b111110001;
assign logo_rueda[22][11] = 9'b101001001;
assign logo_rueda[22][12] = 9'b101001001;
assign logo_rueda[22][13] = 9'b101001000;
assign logo_rueda[22][14] = 9'b110100100;
assign logo_rueda[22][15] = 9'b111111101;
assign logo_rueda[22][16] = 9'b111111110;
assign logo_rueda[22][17] = 9'b111110001;
assign logo_rueda[22][18] = 9'b111111100;
assign logo_rueda[22][19] = 9'b111101100;
assign logo_rueda[22][20] = 9'b111100100;
assign logo_rueda[22][21] = 9'b111101101;
assign logo_rueda[22][22] = 9'b111111110;
assign logo_rueda[22][23] = 9'b111111111;
assign logo_rueda[22][24] = 9'b111101101;
assign logo_rueda[22][25] = 9'b111101000;
assign logo_rueda[22][26] = 9'b111101000;
assign logo_rueda[22][27] = 9'b111101000;
assign logo_rueda[22][28] = 9'b110001000;
assign logo_rueda[22][29] = 9'b100000100;
assign logo_rueda[22][30] = 9'b101001001;
assign logo_rueda[22][31] = 9'b101101000;
assign logo_rueda[22][32] = 9'b101100100;
assign logo_rueda[22][33] = 9'b101100100;
assign logo_rueda[22][34] = 9'b110001000;
assign logo_rueda[22][35] = 9'b101100100;
assign logo_rueda[22][36] = 9'b111111100;
assign logo_rueda[22][37] = 9'b111111100;
assign logo_rueda[22][38] = 9'b111111100;
assign logo_rueda[23][6] = 9'b110101000;
assign logo_rueda[23][7] = 9'b111110100;
assign logo_rueda[23][9] = 9'b110001000;
assign logo_rueda[23][10] = 9'b111111100;
assign logo_rueda[23][11] = 9'b101101101;
assign logo_rueda[23][12] = 9'b101001001;
assign logo_rueda[23][13] = 9'b101001001;
assign logo_rueda[23][14] = 9'b101000100;
assign logo_rueda[23][15] = 9'b111101000;
assign logo_rueda[23][16] = 9'b111111110;
assign logo_rueda[23][17] = 9'b111110001;
assign logo_rueda[23][18] = 9'b111110000;
assign logo_rueda[23][19] = 9'b111101000;
assign logo_rueda[23][20] = 9'b111101101;
assign logo_rueda[23][21] = 9'b111110001;
assign logo_rueda[23][22] = 9'b111101101;
assign logo_rueda[23][23] = 9'b111111101;
assign logo_rueda[23][24] = 9'b111110101;
assign logo_rueda[23][25] = 9'b111110101;
assign logo_rueda[23][26] = 9'b111111111;
assign logo_rueda[23][27] = 9'b111110101;
assign logo_rueda[23][28] = 9'b111101101;
assign logo_rueda[23][29] = 9'b100100100;
assign logo_rueda[23][30] = 9'b100100100;
assign logo_rueda[23][31] = 9'b101001000;
assign logo_rueda[23][32] = 9'b110001000;
assign logo_rueda[23][33] = 9'b101000100;
assign logo_rueda[23][34] = 9'b110001000;
assign logo_rueda[23][35] = 9'b101000100;
assign logo_rueda[23][36] = 9'b110001000;
assign logo_rueda[23][37] = 9'b111111100;
assign logo_rueda[23][38] = 9'b111110100;
assign logo_rueda[24][6] = 9'b101000000;
assign logo_rueda[24][7] = 9'b111110000;
assign logo_rueda[24][8] = 9'b111110001;
assign logo_rueda[24][9] = 9'b100100000;
assign logo_rueda[24][10] = 9'b111110000;
assign logo_rueda[24][11] = 9'b111110001;
assign logo_rueda[24][12] = 9'b101001001;
assign logo_rueda[24][13] = 9'b101001001;
assign logo_rueda[24][14] = 9'b101001001;
assign logo_rueda[24][15] = 9'b101100100;
assign logo_rueda[24][16] = 9'b111110001;
assign logo_rueda[24][17] = 9'b111111101;
assign logo_rueda[24][18] = 9'b111101000;
assign logo_rueda[24][19] = 9'b111101101;
assign logo_rueda[24][20] = 9'b111111110;
assign logo_rueda[24][21] = 9'b111111111;
assign logo_rueda[24][22] = 9'b111110001;
assign logo_rueda[24][23] = 9'b111101101;
assign logo_rueda[24][24] = 9'b111110001;
assign logo_rueda[24][25] = 9'b111110101;
assign logo_rueda[24][26] = 9'b111111111;
assign logo_rueda[24][27] = 9'b111111111;
assign logo_rueda[24][28] = 9'b111111101;
assign logo_rueda[24][29] = 9'b101101000;
assign logo_rueda[24][30] = 9'b100000000;
assign logo_rueda[24][31] = 9'b101001001;
assign logo_rueda[24][32] = 9'b101000100;
assign logo_rueda[24][33] = 9'b110001000;
assign logo_rueda[24][34] = 9'b101000100;
assign logo_rueda[24][35] = 9'b110001000;
assign logo_rueda[24][36] = 9'b100100000;
assign logo_rueda[24][37] = 9'b111110100;
assign logo_rueda[24][38] = 9'b111111100;
assign logo_rueda[24][39] = 9'b110000100;
assign logo_rueda[24][40] = 9'b111101000;
assign logo_rueda[25][7] = 9'b110000100;
assign logo_rueda[25][8] = 9'b111110000;
assign logo_rueda[25][10] = 9'b110000100;
assign logo_rueda[25][11] = 9'b111110100;
assign logo_rueda[25][12] = 9'b110001101;
assign logo_rueda[25][13] = 9'b101001001;
assign logo_rueda[25][14] = 9'b101001101;
assign logo_rueda[25][15] = 9'b101001000;
assign logo_rueda[25][16] = 9'b110000000;
assign logo_rueda[25][17] = 9'b111110001;
assign logo_rueda[25][18] = 9'b110101101;
assign logo_rueda[25][19] = 9'b111110001;
assign logo_rueda[25][20] = 9'b111111111;
assign logo_rueda[25][21] = 9'b111111111;
assign logo_rueda[25][22] = 9'b111110101;
assign logo_rueda[25][23] = 9'b111101000;
assign logo_rueda[25][24] = 9'b111101100;
assign logo_rueda[25][25] = 9'b111101100;
assign logo_rueda[25][26] = 9'b111110001;
assign logo_rueda[25][27] = 9'b111111110;
assign logo_rueda[25][28] = 9'b111111101;
assign logo_rueda[25][29] = 9'b111101100;
assign logo_rueda[25][30] = 9'b100100000;
assign logo_rueda[25][31] = 9'b101001001;
assign logo_rueda[25][32] = 9'b101001001;
assign logo_rueda[25][33] = 9'b101100100;
assign logo_rueda[25][34] = 9'b110001000;
assign logo_rueda[25][35] = 9'b110000100;
assign logo_rueda[25][36] = 9'b101000100;
assign logo_rueda[25][37] = 9'b101100100;
assign logo_rueda[25][38] = 9'b111110100;
assign logo_rueda[25][39] = 9'b110000100;
assign logo_rueda[25][40] = 9'b111101100;
assign logo_rueda[26][7] = 9'b100100000;
assign logo_rueda[26][8] = 9'b111101100;
assign logo_rueda[26][9] = 9'b111110001;
assign logo_rueda[26][10] = 9'b100000000;
assign logo_rueda[26][11] = 9'b111101100;
assign logo_rueda[26][12] = 9'b111110000;
assign logo_rueda[26][13] = 9'b101001001;
assign logo_rueda[26][14] = 9'b101001001;
assign logo_rueda[26][15] = 9'b101001101;
assign logo_rueda[26][16] = 9'b101000100;
assign logo_rueda[26][17] = 9'b110000100;
assign logo_rueda[26][18] = 9'b111110001;
assign logo_rueda[26][19] = 9'b110110001;
assign logo_rueda[26][20] = 9'b111111111;
assign logo_rueda[26][21] = 9'b111111111;
assign logo_rueda[26][22] = 9'b111101100;
assign logo_rueda[26][23] = 9'b111101000;
assign logo_rueda[26][24] = 9'b111110101;
assign logo_rueda[26][25] = 9'b111110001;
assign logo_rueda[26][26] = 9'b111101000;
assign logo_rueda[26][27] = 9'b111110001;
assign logo_rueda[26][28] = 9'b111110001;
assign logo_rueda[26][29] = 9'b111101101;
assign logo_rueda[26][30] = 9'b101000100;
assign logo_rueda[26][31] = 9'b100100100;
assign logo_rueda[26][32] = 9'b101001101;
assign logo_rueda[26][33] = 9'b100100100;
assign logo_rueda[26][34] = 9'b110001000;
assign logo_rueda[26][35] = 9'b101100100;
assign logo_rueda[26][36] = 9'b101100100;
assign logo_rueda[26][37] = 9'b100100000;
assign logo_rueda[26][38] = 9'b111101100;
assign logo_rueda[26][39] = 9'b110001000;
assign logo_rueda[26][40] = 9'b110101000;
assign logo_rueda[27][8] = 9'b101000000;
assign logo_rueda[27][9] = 9'b111101100;
assign logo_rueda[27][11] = 9'b101100000;
assign logo_rueda[27][12] = 9'b111110100;
assign logo_rueda[27][13] = 9'b110001101;
assign logo_rueda[27][14] = 9'b101001001;
assign logo_rueda[27][15] = 9'b101001101;
assign logo_rueda[27][16] = 9'b101001001;
assign logo_rueda[27][17] = 9'b100100000;
assign logo_rueda[27][18] = 9'b110100100;
assign logo_rueda[27][19] = 9'b111101100;
assign logo_rueda[27][20] = 9'b111110101;
assign logo_rueda[27][21] = 9'b111110001;
assign logo_rueda[27][22] = 9'b111101100;
assign logo_rueda[27][23] = 9'b111101100;
assign logo_rueda[27][24] = 9'b111110001;
assign logo_rueda[27][25] = 9'b111111111;
assign logo_rueda[27][26] = 9'b111101100;
assign logo_rueda[27][27] = 9'b111110000;
assign logo_rueda[27][28] = 9'b111111100;
assign logo_rueda[27][29] = 9'b111110101;
assign logo_rueda[27][30] = 9'b101101000;
assign logo_rueda[27][31] = 9'b100000000;
assign logo_rueda[27][32] = 9'b101001001;
assign logo_rueda[27][33] = 9'b101001001;
assign logo_rueda[27][34] = 9'b101000100;
assign logo_rueda[27][35] = 9'b110001000;
assign logo_rueda[27][36] = 9'b101100100;
assign logo_rueda[27][37] = 9'b110000100;
assign logo_rueda[27][38] = 9'b111110000;
assign logo_rueda[27][39] = 9'b110001000;
assign logo_rueda[27][40] = 9'b110001000;
assign logo_rueda[28][9] = 9'b101100100;
assign logo_rueda[28][10] = 9'b111101100;
assign logo_rueda[28][12] = 9'b110001000;
assign logo_rueda[28][13] = 9'b111110100;
assign logo_rueda[28][14] = 9'b101101001;
assign logo_rueda[28][15] = 9'b101001001;
assign logo_rueda[28][16] = 9'b101101101;
assign logo_rueda[28][17] = 9'b100100100;
assign logo_rueda[28][18] = 9'b100100100;
assign logo_rueda[28][19] = 9'b110100100;
assign logo_rueda[28][20] = 9'b111101000;
assign logo_rueda[28][21] = 9'b111101100;
assign logo_rueda[28][22] = 9'b111111100;
assign logo_rueda[28][23] = 9'b111111100;
assign logo_rueda[28][24] = 9'b111110000;
assign logo_rueda[28][25] = 9'b111111110;
assign logo_rueda[28][26] = 9'b111111110;
assign logo_rueda[28][27] = 9'b111101100;
assign logo_rueda[28][28] = 9'b111111100;
assign logo_rueda[28][29] = 9'b111111100;
assign logo_rueda[28][30] = 9'b110001100;
assign logo_rueda[28][31] = 9'b100000000;
assign logo_rueda[28][32] = 9'b101101101;
assign logo_rueda[28][33] = 9'b110110110;
assign logo_rueda[28][34] = 9'b101001000;
assign logo_rueda[28][35] = 9'b110001000;
assign logo_rueda[28][36] = 9'b110001000;
assign logo_rueda[28][37] = 9'b100100000;
assign logo_rueda[28][38] = 9'b111101100;
assign logo_rueda[28][39] = 9'b110101100;
assign logo_rueda[28][40] = 9'b110000100;
assign logo_rueda[28][41] = 9'b111110001;
assign logo_rueda[29][10] = 9'b101100100;
assign logo_rueda[29][11] = 9'b111101100;
assign logo_rueda[29][12] = 9'b100100000;
assign logo_rueda[29][13] = 9'b111101100;
assign logo_rueda[29][14] = 9'b111110000;
assign logo_rueda[29][15] = 9'b101001001;
assign logo_rueda[29][16] = 9'b101001101;
assign logo_rueda[29][17] = 9'b101001001;
assign logo_rueda[29][18] = 9'b100101000;
assign logo_rueda[29][19] = 9'b100100100;
assign logo_rueda[29][20] = 9'b110000000;
assign logo_rueda[29][21] = 9'b111101000;
assign logo_rueda[29][22] = 9'b111111100;
assign logo_rueda[29][23] = 9'b111111100;
assign logo_rueda[29][24] = 9'b111110100;
assign logo_rueda[29][25] = 9'b111110001;
assign logo_rueda[29][26] = 9'b111111111;
assign logo_rueda[29][27] = 9'b111110001;
assign logo_rueda[29][28] = 9'b111110100;
assign logo_rueda[29][29] = 9'b111111100;
assign logo_rueda[29][30] = 9'b110101000;
assign logo_rueda[29][31] = 9'b100000000;
assign logo_rueda[29][32] = 9'b101101101;
assign logo_rueda[29][33] = 9'b110010001;
assign logo_rueda[29][34] = 9'b101101101;
assign logo_rueda[29][35] = 9'b101000100;
assign logo_rueda[29][36] = 9'b110101100;
assign logo_rueda[29][37] = 9'b100000000;
assign logo_rueda[29][38] = 9'b101100100;
assign logo_rueda[29][39] = 9'b111110000;
assign logo_rueda[29][40] = 9'b101100100;
assign logo_rueda[29][41] = 9'b111101100;
assign logo_rueda[30][11] = 9'b110000100;
assign logo_rueda[30][12] = 9'b111101000;
assign logo_rueda[30][13] = 9'b101000000;
assign logo_rueda[30][14] = 9'b111110000;
assign logo_rueda[30][15] = 9'b110001100;
assign logo_rueda[30][16] = 9'b101001001;
assign logo_rueda[30][17] = 9'b101001001;
assign logo_rueda[30][18] = 9'b101101001;
assign logo_rueda[30][19] = 9'b101001001;
assign logo_rueda[30][20] = 9'b100100100;
assign logo_rueda[30][21] = 9'b101100100;
assign logo_rueda[30][22] = 9'b111100100;
assign logo_rueda[30][23] = 9'b111101100;
assign logo_rueda[30][24] = 9'b111110000;
assign logo_rueda[30][25] = 9'b111110000;
assign logo_rueda[30][26] = 9'b111110101;
assign logo_rueda[30][27] = 9'b111111101;
assign logo_rueda[30][28] = 9'b111101100;
assign logo_rueda[30][29] = 9'b111111100;
assign logo_rueda[30][30] = 9'b110000100;
assign logo_rueda[30][31] = 9'b100000000;
assign logo_rueda[30][32] = 9'b101101101;
assign logo_rueda[30][33] = 9'b110010010;
assign logo_rueda[30][34] = 9'b101101101;
assign logo_rueda[30][35] = 9'b100100000;
assign logo_rueda[30][36] = 9'b110101000;
assign logo_rueda[30][37] = 9'b100100100;
assign logo_rueda[30][38] = 9'b100100000;
assign logo_rueda[30][39] = 9'b111110000;
assign logo_rueda[30][40] = 9'b110001000;
assign logo_rueda[30][41] = 9'b110101100;
assign logo_rueda[31][14] = 9'b101100000;
assign logo_rueda[31][15] = 9'b111110000;
assign logo_rueda[31][16] = 9'b101101000;
assign logo_rueda[31][17] = 9'b100100100;
assign logo_rueda[31][18] = 9'b101101101;
assign logo_rueda[31][19] = 9'b101101101;
assign logo_rueda[31][20] = 9'b101001001;
assign logo_rueda[31][21] = 9'b101001001;
assign logo_rueda[31][22] = 9'b101101000;
assign logo_rueda[31][23] = 9'b110000100;
assign logo_rueda[31][24] = 9'b111100000;
assign logo_rueda[31][25] = 9'b111100100;
assign logo_rueda[31][26] = 9'b111101100;
assign logo_rueda[31][27] = 9'b111110001;
assign logo_rueda[31][28] = 9'b111101100;
assign logo_rueda[31][29] = 9'b111101000;
assign logo_rueda[31][30] = 9'b101000100;
assign logo_rueda[31][31] = 9'b100000100;
assign logo_rueda[31][32] = 9'b101101101;
assign logo_rueda[31][33] = 9'b110010001;
assign logo_rueda[31][34] = 9'b101101101;
assign logo_rueda[31][35] = 9'b100000000;
assign logo_rueda[31][36] = 9'b101100100;
assign logo_rueda[31][37] = 9'b101101000;
assign logo_rueda[31][38] = 9'b100000000;
assign logo_rueda[31][39] = 9'b111101100;
assign logo_rueda[31][40] = 9'b110110000;
assign logo_rueda[31][41] = 9'b110000100;
assign logo_rueda[31][42] = 9'b111110000;
assign logo_rueda[32][15] = 9'b101100100;
assign logo_rueda[32][16] = 9'b111110000;
assign logo_rueda[32][17] = 9'b101000100;
assign logo_rueda[32][18] = 9'b101001001;
assign logo_rueda[32][19] = 9'b110010001;
assign logo_rueda[32][20] = 9'b110010010;
assign logo_rueda[32][21] = 9'b110010010;
assign logo_rueda[32][22] = 9'b101101101;
assign logo_rueda[32][23] = 9'b101101101;
assign logo_rueda[32][24] = 9'b101101000;
assign logo_rueda[32][25] = 9'b110000100;
assign logo_rueda[32][26] = 9'b110100100;
assign logo_rueda[32][27] = 9'b111100100;
assign logo_rueda[32][28] = 9'b110100100;
assign logo_rueda[32][29] = 9'b101100100;
assign logo_rueda[32][30] = 9'b100100100;
assign logo_rueda[32][31] = 9'b101001001;
assign logo_rueda[32][32] = 9'b101101101;
assign logo_rueda[32][33] = 9'b110010001;
assign logo_rueda[32][34] = 9'b101101101;
assign logo_rueda[32][35] = 9'b100100100;
assign logo_rueda[32][36] = 9'b101000100;
assign logo_rueda[32][37] = 9'b110101100;
assign logo_rueda[32][38] = 9'b100000000;
assign logo_rueda[32][39] = 9'b110001000;
assign logo_rueda[32][40] = 9'b111110100;
assign logo_rueda[32][41] = 9'b110000100;
assign logo_rueda[32][42] = 9'b111110000;
assign logo_rueda[32][43] = 9'b111101101;
assign logo_rueda[33][16] = 9'b101100100;
assign logo_rueda[33][17] = 9'b111110000;
assign logo_rueda[33][18] = 9'b101000100;
assign logo_rueda[33][19] = 9'b100100100;
assign logo_rueda[33][20] = 9'b101101101;
assign logo_rueda[33][21] = 9'b111111111;
assign logo_rueda[33][22] = 9'b110010001;
assign logo_rueda[33][23] = 9'b110010001;
assign logo_rueda[33][24] = 9'b110010001;
assign logo_rueda[33][25] = 9'b101001001;
assign logo_rueda[33][26] = 9'b101101001;
assign logo_rueda[33][27] = 9'b101001000;
assign logo_rueda[33][28] = 9'b101001000;
assign logo_rueda[33][29] = 9'b100101000;
assign logo_rueda[33][30] = 9'b101001001;
assign logo_rueda[33][31] = 9'b110010001;
assign logo_rueda[33][32] = 9'b101101101;
assign logo_rueda[33][33] = 9'b110010001;
assign logo_rueda[33][34] = 9'b101001000;
assign logo_rueda[33][35] = 9'b100100100;
assign logo_rueda[33][36] = 9'b101000100;
assign logo_rueda[33][37] = 9'b111101100;
assign logo_rueda[33][38] = 9'b100000000;
assign logo_rueda[33][39] = 9'b101100100;
assign logo_rueda[33][40] = 9'b110101000;
assign logo_rueda[33][41] = 9'b111101100;
assign logo_rueda[33][42] = 9'b111101100;
assign logo_rueda[33][43] = 9'b111110000;
assign logo_rueda[34][17] = 9'b101100100;
assign logo_rueda[34][18] = 9'b111101100;
assign logo_rueda[34][19] = 9'b100100100;
assign logo_rueda[34][20] = 9'b100000000;
assign logo_rueda[34][21] = 9'b101101101;
assign logo_rueda[34][22] = 9'b110010010;
assign logo_rueda[34][23] = 9'b101001001;
assign logo_rueda[34][24] = 9'b101101101;
assign logo_rueda[34][25] = 9'b110110110;
assign logo_rueda[34][26] = 9'b101001001;
assign logo_rueda[34][27] = 9'b101101101;
assign logo_rueda[34][28] = 9'b101101101;
assign logo_rueda[34][29] = 9'b110010001;
assign logo_rueda[34][30] = 9'b110010010;
assign logo_rueda[34][31] = 9'b101001001;
assign logo_rueda[34][32] = 9'b110010001;
assign logo_rueda[34][33] = 9'b101101101;
assign logo_rueda[34][34] = 9'b101001001;
assign logo_rueda[34][35] = 9'b100100100;
assign logo_rueda[34][36] = 9'b101000000;
assign logo_rueda[34][37] = 9'b111110000;
assign logo_rueda[34][38] = 9'b100000000;
assign logo_rueda[34][39] = 9'b100100000;
assign logo_rueda[34][40] = 9'b101000000;
assign logo_rueda[34][41] = 9'b111110000;
assign logo_rueda[34][42] = 9'b111111100;
assign logo_rueda[34][43] = 9'b111110000;
assign logo_rueda[35][17] = 9'b100000000;
assign logo_rueda[35][18] = 9'b101100100;
assign logo_rueda[35][19] = 9'b111101100;
assign logo_rueda[35][20] = 9'b101000100;
assign logo_rueda[35][21] = 9'b100100100;
assign logo_rueda[35][22] = 9'b101101101;
assign logo_rueda[35][23] = 9'b101101101;
assign logo_rueda[35][24] = 9'b101101101;
assign logo_rueda[35][25] = 9'b101001001;
assign logo_rueda[35][26] = 9'b100100100;
assign logo_rueda[35][27] = 9'b101101101;
assign logo_rueda[35][28] = 9'b101101101;
assign logo_rueda[35][29] = 9'b101001001;
assign logo_rueda[35][30] = 9'b101101101;
assign logo_rueda[35][31] = 9'b101001001;
assign logo_rueda[35][32] = 9'b101001000;
assign logo_rueda[35][33] = 9'b100100100;
assign logo_rueda[35][34] = 9'b100100100;
assign logo_rueda[35][35] = 9'b100100100;
assign logo_rueda[35][36] = 9'b101000100;
assign logo_rueda[35][37] = 9'b111110000;
assign logo_rueda[35][38] = 9'b100100000;
assign logo_rueda[35][39] = 9'b100000000;
assign logo_rueda[35][40] = 9'b100000000;
assign logo_rueda[35][41] = 9'b110001000;
assign logo_rueda[35][42] = 9'b111111100;
assign logo_rueda[35][43] = 9'b111110100;
assign logo_rueda[35][44] = 9'b111101101;
assign logo_rueda[36][18] = 9'b100000000;
assign logo_rueda[36][19] = 9'b101000000;
assign logo_rueda[36][20] = 9'b111101000;
assign logo_rueda[36][21] = 9'b101101000;
assign logo_rueda[36][22] = 9'b100000000;
assign logo_rueda[36][23] = 9'b100101000;
assign logo_rueda[36][24] = 9'b101101101;
assign logo_rueda[36][25] = 9'b100000100;
assign logo_rueda[36][26] = 9'b101101101;
assign logo_rueda[36][27] = 9'b110010001;
assign logo_rueda[36][28] = 9'b101001001;
assign logo_rueda[36][29] = 9'b101001001;
assign logo_rueda[36][30] = 9'b101001001;
assign logo_rueda[36][31] = 9'b101001000;
assign logo_rueda[36][32] = 9'b101001000;
assign logo_rueda[36][33] = 9'b100100100;
assign logo_rueda[36][34] = 9'b100000000;
assign logo_rueda[36][35] = 9'b100000000;
assign logo_rueda[36][36] = 9'b110001000;
assign logo_rueda[36][37] = 9'b111110000;
assign logo_rueda[36][38] = 9'b100000000;
assign logo_rueda[36][39] = 9'b100000000;
assign logo_rueda[36][40] = 9'b100000000;
assign logo_rueda[36][41] = 9'b101100100;
assign logo_rueda[36][42] = 9'b111110000;
assign logo_rueda[36][43] = 9'b111110000;
assign logo_rueda[36][44] = 9'b111110000;
assign logo_rueda[37][18] = 9'b111101000;
assign logo_rueda[37][19] = 9'b101000100;
assign logo_rueda[37][20] = 9'b100000000;
assign logo_rueda[37][21] = 9'b110001000;
assign logo_rueda[37][22] = 9'b110001000;
assign logo_rueda[37][23] = 9'b100100000;
assign logo_rueda[37][24] = 9'b100000100;
assign logo_rueda[37][25] = 9'b100100100;
assign logo_rueda[37][26] = 9'b100100100;
assign logo_rueda[37][27] = 9'b101001001;
assign logo_rueda[37][28] = 9'b101101101;
assign logo_rueda[37][29] = 9'b100100100;
assign logo_rueda[37][30] = 9'b100100100;
assign logo_rueda[37][31] = 9'b100000000;
assign logo_rueda[37][32] = 9'b100100100;
assign logo_rueda[37][33] = 9'b100100100;
assign logo_rueda[37][34] = 9'b100000000;
assign logo_rueda[37][35] = 9'b100100000;
assign logo_rueda[37][36] = 9'b111110000;
assign logo_rueda[37][37] = 9'b111110000;
assign logo_rueda[37][38] = 9'b100000000;
assign logo_rueda[37][39] = 9'b100000000;
assign logo_rueda[37][40] = 9'b100000000;
assign logo_rueda[37][41] = 9'b101000100;
assign logo_rueda[37][42] = 9'b111110000;
assign logo_rueda[37][43] = 9'b111110000;
assign logo_rueda[37][44] = 9'b111110000;
assign logo_rueda[38][18] = 9'b101100100;
assign logo_rueda[38][19] = 9'b111101000;
assign logo_rueda[38][20] = 9'b110001000;
assign logo_rueda[38][21] = 9'b100000000;
assign logo_rueda[38][22] = 9'b101000000;
assign logo_rueda[38][23] = 9'b101100100;
assign logo_rueda[38][24] = 9'b100000000;
assign logo_rueda[38][25] = 9'b100100100;
assign logo_rueda[38][26] = 9'b100000000;
assign logo_rueda[38][27] = 9'b100000000;
assign logo_rueda[38][28] = 9'b100100100;
assign logo_rueda[38][29] = 9'b100000000;
assign logo_rueda[38][30] = 9'b100000000;
assign logo_rueda[38][31] = 9'b100000000;
assign logo_rueda[38][32] = 9'b100000000;
assign logo_rueda[38][33] = 9'b100000000;
assign logo_rueda[38][34] = 9'b100000000;
assign logo_rueda[38][35] = 9'b110001000;
assign logo_rueda[38][36] = 9'b111110100;
assign logo_rueda[38][37] = 9'b101000100;
assign logo_rueda[38][38] = 9'b100000000;
assign logo_rueda[38][39] = 9'b100000000;
assign logo_rueda[38][40] = 9'b100000000;
assign logo_rueda[38][41] = 9'b101100100;
assign logo_rueda[38][42] = 9'b111110000;
assign logo_rueda[38][43] = 9'b111101100;
assign logo_rueda[38][44] = 9'b111110000;
assign logo_rueda[39][19] = 9'b101000000;
assign logo_rueda[39][20] = 9'b111101100;
assign logo_rueda[39][21] = 9'b111110000;
assign logo_rueda[39][22] = 9'b101000100;
assign logo_rueda[39][23] = 9'b100000000;
assign logo_rueda[39][24] = 9'b100000000;
assign logo_rueda[39][25] = 9'b100000000;
assign logo_rueda[39][26] = 9'b100000000;
assign logo_rueda[39][27] = 9'b100000000;
assign logo_rueda[39][28] = 9'b100000000;
assign logo_rueda[39][29] = 9'b100100100;
assign logo_rueda[39][30] = 9'b100000000;
assign logo_rueda[39][31] = 9'b100000000;
assign logo_rueda[39][32] = 9'b100000000;
assign logo_rueda[39][33] = 9'b100100100;
assign logo_rueda[39][34] = 9'b100000100;
assign logo_rueda[39][35] = 9'b101000000;
assign logo_rueda[39][36] = 9'b101000000;
assign logo_rueda[39][37] = 9'b101100100;
assign logo_rueda[39][38] = 9'b100000000;
assign logo_rueda[39][39] = 9'b100000000;
assign logo_rueda[39][40] = 9'b100000000;
assign logo_rueda[39][41] = 9'b110001000;
assign logo_rueda[39][42] = 9'b111110000;
assign logo_rueda[39][43] = 9'b111101100;
assign logo_rueda[39][44] = 9'b111110000;
assign logo_rueda[40][20] = 9'b101000000;
assign logo_rueda[40][21] = 9'b110101000;
assign logo_rueda[40][22] = 9'b111110100;
assign logo_rueda[40][23] = 9'b111110000;
assign logo_rueda[40][24] = 9'b101100100;
assign logo_rueda[40][25] = 9'b100100000;
assign logo_rueda[40][26] = 9'b100000000;
assign logo_rueda[40][27] = 9'b100000000;
assign logo_rueda[40][28] = 9'b100000000;
assign logo_rueda[40][29] = 9'b100000000;
assign logo_rueda[40][30] = 9'b100000000;
assign logo_rueda[40][31] = 9'b100000000;
assign logo_rueda[40][32] = 9'b100000000;
assign logo_rueda[40][33] = 9'b100000000;
assign logo_rueda[40][34] = 9'b100000000;
assign logo_rueda[40][35] = 9'b100100000;
assign logo_rueda[40][36] = 9'b110101100;
assign logo_rueda[40][37] = 9'b110101100;
assign logo_rueda[40][38] = 9'b100000000;
assign logo_rueda[40][39] = 9'b100000000;
assign logo_rueda[40][40] = 9'b100000000;
assign logo_rueda[40][41] = 9'b111101100;
assign logo_rueda[40][42] = 9'b111101100;
assign logo_rueda[40][43] = 9'b111101100;
assign logo_rueda[40][44] = 9'b111110000;
assign logo_rueda[41][22] = 9'b110000100;
assign logo_rueda[41][23] = 9'b111110000;
assign logo_rueda[41][24] = 9'b111111100;
assign logo_rueda[41][25] = 9'b111110100;
assign logo_rueda[41][26] = 9'b110101100;
assign logo_rueda[41][27] = 9'b101101000;
assign logo_rueda[41][28] = 9'b101000100;
assign logo_rueda[41][29] = 9'b100100000;
assign logo_rueda[41][30] = 9'b100100000;
assign logo_rueda[41][31] = 9'b100100000;
assign logo_rueda[41][32] = 9'b101000100;
assign logo_rueda[41][33] = 9'b101100100;
assign logo_rueda[41][34] = 9'b110101100;
assign logo_rueda[41][35] = 9'b111110100;
assign logo_rueda[41][36] = 9'b111110000;
assign logo_rueda[41][37] = 9'b100100000;
assign logo_rueda[41][38] = 9'b100000000;
assign logo_rueda[41][39] = 9'b100000000;
assign logo_rueda[41][40] = 9'b110001000;
assign logo_rueda[41][41] = 9'b111110000;
assign logo_rueda[41][42] = 9'b111101100;
assign logo_rueda[41][43] = 9'b111101100;
assign logo_rueda[41][44] = 9'b111110000;
assign logo_rueda[42][23] = 9'b101100000;
assign logo_rueda[42][24] = 9'b110101000;
assign logo_rueda[42][25] = 9'b111110000;
assign logo_rueda[42][26] = 9'b111110100;
assign logo_rueda[42][27] = 9'b111110000;
assign logo_rueda[42][28] = 9'b111110000;
assign logo_rueda[42][29] = 9'b111110000;
assign logo_rueda[42][30] = 9'b111110000;
assign logo_rueda[42][31] = 9'b111110000;
assign logo_rueda[42][32] = 9'b111110000;
assign logo_rueda[42][33] = 9'b111110000;
assign logo_rueda[42][34] = 9'b111110000;
assign logo_rueda[42][35] = 9'b111110000;
assign logo_rueda[42][36] = 9'b100000000;
assign logo_rueda[42][37] = 9'b100000000;
assign logo_rueda[42][38] = 9'b100000000;
assign logo_rueda[42][39] = 9'b110001000;
assign logo_rueda[42][40] = 9'b111110000;
assign logo_rueda[42][41] = 9'b111101100;
assign logo_rueda[42][42] = 9'b111101000;
assign logo_rueda[42][43] = 9'b111101000;
assign logo_rueda[42][44] = 9'b111110000;
assign logo_rueda[43][25] = 9'b101100000;
assign logo_rueda[43][26] = 9'b110101000;
assign logo_rueda[43][27] = 9'b111101100;
assign logo_rueda[43][28] = 9'b111101100;
assign logo_rueda[43][29] = 9'b111101100;
assign logo_rueda[43][30] = 9'b111101100;
assign logo_rueda[43][31] = 9'b111101000;
assign logo_rueda[43][32] = 9'b111100100;
assign logo_rueda[43][33] = 9'b111100100;
assign logo_rueda[43][34] = 9'b111101000;
assign logo_rueda[43][35] = 9'b111110000;
assign logo_rueda[43][36] = 9'b110001000;
assign logo_rueda[43][37] = 9'b110001100;
assign logo_rueda[43][38] = 9'b111110000;
assign logo_rueda[43][39] = 9'b111110100;
assign logo_rueda[43][40] = 9'b111101100;
assign logo_rueda[43][41] = 9'b111101100;
assign logo_rueda[43][42] = 9'b111101100;
assign logo_rueda[43][43] = 9'b111101100;
assign logo_rueda[43][44] = 9'b111110000;
assign logo_rueda[44][27] = 9'b101100000;
assign logo_rueda[44][28] = 9'b110000100;
assign logo_rueda[44][29] = 9'b110101000;
assign logo_rueda[44][30] = 9'b111101100;
assign logo_rueda[44][31] = 9'b111101100;
assign logo_rueda[44][32] = 9'b111101100;
assign logo_rueda[44][33] = 9'b111110000;
assign logo_rueda[44][34] = 9'b111110000;
assign logo_rueda[44][35] = 9'b111110000;
assign logo_rueda[44][36] = 9'b111110100;
assign logo_rueda[44][37] = 9'b111110100;
assign logo_rueda[44][38] = 9'b111110000;
assign logo_rueda[44][39] = 9'b111110000;
assign logo_rueda[44][40] = 9'b111110100;
assign logo_rueda[44][41] = 9'b111101100;
assign logo_rueda[44][42] = 9'b111101000;
assign logo_rueda[44][43] = 9'b111101100;
assign logo_rueda[44][44] = 9'b111110000;
assign logo_rueda[45][30] = 9'b101100000;
assign logo_rueda[45][31] = 9'b110000100;
assign logo_rueda[45][32] = 9'b110001000;
assign logo_rueda[45][33] = 9'b110101000;
assign logo_rueda[45][34] = 9'b110101000;
assign logo_rueda[45][35] = 9'b110100100;
assign logo_rueda[45][36] = 9'b110100100;
assign logo_rueda[45][37] = 9'b110000000;
assign logo_rueda[45][38] = 9'b110000000;
assign logo_rueda[45][39] = 9'b101100100;
assign logo_rueda[45][40] = 9'b111101100;
assign logo_rueda[45][41] = 9'b111110000;
assign logo_rueda[45][42] = 9'b111101100;
assign logo_rueda[45][43] = 9'b111110000;
assign logo_rueda[45][44] = 9'b111101100;
assign logo_rueda[46][40] = 9'b110101000;
assign logo_rueda[46][41] = 9'b111110000;
assign logo_rueda[46][42] = 9'b111110100;
assign logo_rueda[46][43] = 9'b111101100;
assign logo_rueda[47][32] = 9'b111101000;
assign logo_rueda[47][38] = 9'b111101100;
assign logo_rueda[47][39] = 9'b111110000;
assign logo_rueda[47][40] = 9'b111111100;
assign logo_rueda[47][41] = 9'b111111100;
assign logo_rueda[47][42] = 9'b111110000;
assign logo_rueda[48][32] = 9'b110000100;
assign logo_rueda[48][33] = 9'b110101000;
assign logo_rueda[48][34] = 9'b111101000;
assign logo_rueda[48][35] = 9'b111101100;
assign logo_rueda[48][36] = 9'b111101100;
assign logo_rueda[48][37] = 9'b111110000;
assign logo_rueda[48][38] = 9'b111110100;
assign logo_rueda[48][39] = 9'b111110100;
assign logo_rueda[48][40] = 9'b111110000;
assign logo_rueda[48][41] = 9'b111101000;
assign logo_rueda[49][35] = 9'b110000100;
assign logo_rueda[49][36] = 9'b110000100;
assign logo_rueda[49][37] = 9'b110101000;
assign logo_rueda[49][38] = 9'b111101000;
//Total de Lineas = 1479
endmodule

