`timescale 1ns / 1ps
module racing (
input enable,
input clock,
input [9:0] posx, posy,
input [9:0] hcount,
input [9:0] vcount,
output reg[2:0] red,
output reg[2:0] green,
output reg[1:0] blue,
output reg data);

always @(posedge clock)
begin
	if(enable)
	begin
		if(hcount >= posx & hcount < posx + RESOLUCION_X & vcount >= posy & vcount < posy + RESOLUCION_Y)
		begin
			if (racing[vcount - posy][hcount - posx][8] == 1'b1)
			begin
				red   <= racing[vcount- posy][hcount- posx][7:5];
				green <= racing[vcount- posy][hcount- posx][4:2];
            blue 	<= racing[vcount- posy][hcount- posx][1:0];
				data  <= 1'b1;
			end
			else
				data <= 0;
			end
		else
		data <= 0;
	end
end

parameter RESOLUCION_X = 25;
parameter RESOLUCION_Y = 50;
wire [8:0] racing[RESOLUCION_Y - 1'b1 : 0][RESOLUCION_X - 1'b1 : 0];
assign racing[2][11] = 9'b100000100;
assign racing[2][12] = 9'b100100100;
assign racing[2][13] = 9'b100100100;
assign racing[2][14] = 9'b100100100;
assign racing[2][15] = 9'b100000100;
assign racing[3][8] = 9'b100000000;
assign racing[3][9] = 9'b100100101;
assign racing[3][10] = 9'b100101001;
assign racing[3][11] = 9'b100101001;
assign racing[3][12] = 9'b100101001;
assign racing[3][13] = 9'b100101001;
assign racing[3][14] = 9'b100101001;
assign racing[3][15] = 9'b100101001;
assign racing[3][16] = 9'b100101001;
assign racing[3][17] = 9'b100100100;
assign racing[4][7] = 9'b100100100;
assign racing[4][8] = 9'b100101001;
assign racing[4][9] = 9'b100101001;
assign racing[4][10] = 9'b100101001;
assign racing[4][11] = 9'b100101001;
assign racing[4][12] = 9'b100101001;
assign racing[4][13] = 9'b100101001;
assign racing[4][14] = 9'b100101001;
assign racing[4][15] = 9'b100101001;
assign racing[4][16] = 9'b100101001;
assign racing[4][17] = 9'b100101001;
assign racing[4][18] = 9'b100101001;
assign racing[5][6] = 9'b100100100;
assign racing[5][7] = 9'b100101001;
assign racing[5][8] = 9'b100101001;
assign racing[5][9] = 9'b100101001;
assign racing[5][10] = 9'b100101001;
assign racing[5][11] = 9'b100101001;
assign racing[5][12] = 9'b100101001;
assign racing[5][13] = 9'b100101001;
assign racing[5][14] = 9'b100101001;
assign racing[5][15] = 9'b100101001;
assign racing[5][16] = 9'b100101001;
assign racing[5][17] = 9'b100101001;
assign racing[5][18] = 9'b100101001;
assign racing[5][19] = 9'b100101001;
assign racing[6][5] = 9'b100000000;
assign racing[6][6] = 9'b100101001;
assign racing[6][7] = 9'b101001001;
assign racing[6][8] = 9'b100101001;
assign racing[6][9] = 9'b100101001;
assign racing[6][10] = 9'b100100101;
assign racing[6][11] = 9'b100100100;
assign racing[6][12] = 9'b100100100;
assign racing[6][13] = 9'b100100100;
assign racing[6][14] = 9'b100100100;
assign racing[6][15] = 9'b100100100;
assign racing[6][16] = 9'b100101001;
assign racing[6][17] = 9'b100101001;
assign racing[6][18] = 9'b100101001;
assign racing[6][19] = 9'b101001001;
assign racing[6][20] = 9'b100100101;
assign racing[7][5] = 9'b100100100;
assign racing[7][6] = 9'b101001001;
assign racing[7][7] = 9'b101001001;
assign racing[7][8] = 9'b100101001;
assign racing[7][9] = 9'b100100101;
assign racing[7][10] = 9'b100000000;
assign racing[7][11] = 9'b100000000;
assign racing[7][12] = 9'b100000000;
assign racing[7][13] = 9'b100000000;
assign racing[7][14] = 9'b100000000;
assign racing[7][15] = 9'b100000000;
assign racing[7][16] = 9'b100100100;
assign racing[7][17] = 9'b100101001;
assign racing[7][18] = 9'b100101001;
assign racing[7][19] = 9'b101001001;
assign racing[7][20] = 9'b100101001;
assign racing[8][5] = 9'b100100101;
assign racing[8][6] = 9'b101001001;
assign racing[8][7] = 9'b101001001;
assign racing[8][8] = 9'b100101001;
assign racing[8][9] = 9'b100100100;
assign racing[8][10] = 9'b100000000;
assign racing[8][11] = 9'b100000000;
assign racing[8][12] = 9'b100000000;
assign racing[8][13] = 9'b100000000;
assign racing[8][14] = 9'b100000000;
assign racing[8][15] = 9'b100000000;
assign racing[8][16] = 9'b100000000;
assign racing[8][17] = 9'b100100101;
assign racing[8][18] = 9'b100101001;
assign racing[8][19] = 9'b101001001;
assign racing[8][20] = 9'b101001001;
assign racing[8][21] = 9'b100100101;
assign racing[9][4] = 9'b100000000;
assign racing[9][5] = 9'b100101001;
assign racing[9][6] = 9'b101001001;
assign racing[9][7] = 9'b101001001;
assign racing[9][8] = 9'b100101001;
assign racing[9][9] = 9'b100100100;
assign racing[9][10] = 9'b100000000;
assign racing[9][11] = 9'b100000000;
assign racing[9][12] = 9'b100000000;
assign racing[9][13] = 9'b100000000;
assign racing[9][14] = 9'b100000000;
assign racing[9][15] = 9'b100000000;
assign racing[9][16] = 9'b100000000;
assign racing[9][17] = 9'b100100100;
assign racing[9][18] = 9'b100101001;
assign racing[9][19] = 9'b101001001;
assign racing[9][20] = 9'b101001001;
assign racing[9][21] = 9'b100101001;
assign racing[10][4] = 9'b100100100;
assign racing[10][5] = 9'b101001001;
assign racing[10][6] = 9'b101001001;
assign racing[10][7] = 9'b101001001;
assign racing[10][8] = 9'b100100101;
assign racing[10][9] = 9'b100000000;
assign racing[10][10] = 9'b100000000;
assign racing[10][11] = 9'b100000000;
assign racing[10][12] = 9'b100000000;
assign racing[10][13] = 9'b100000000;
assign racing[10][14] = 9'b100000000;
assign racing[10][15] = 9'b100000000;
assign racing[10][16] = 9'b100000000;
assign racing[10][17] = 9'b100100100;
assign racing[10][18] = 9'b100101001;
assign racing[10][19] = 9'b101001001;
assign racing[10][20] = 9'b101001001;
assign racing[10][21] = 9'b100101001;
assign racing[11][4] = 9'b100100100;
assign racing[11][5] = 9'b101001001;
assign racing[11][6] = 9'b101001001;
assign racing[11][7] = 9'b101001001;
assign racing[11][8] = 9'b100100100;
assign racing[11][9] = 9'b100000000;
assign racing[11][10] = 9'b100000000;
assign racing[11][11] = 9'b100000000;
assign racing[11][12] = 9'b100000000;
assign racing[11][13] = 9'b100000000;
assign racing[11][14] = 9'b100000000;
assign racing[11][15] = 9'b100000000;
assign racing[11][16] = 9'b100000000;
assign racing[11][17] = 9'b100100100;
assign racing[11][18] = 9'b100101001;
assign racing[11][19] = 9'b101001001;
assign racing[11][20] = 9'b101001001;
assign racing[11][21] = 9'b100101001;
assign racing[12][4] = 9'b100100100;
assign racing[12][5] = 9'b101001001;
assign racing[12][6] = 9'b101001001;
assign racing[12][7] = 9'b100101001;
assign racing[12][8] = 9'b100100100;
assign racing[12][9] = 9'b100000000;
assign racing[12][10] = 9'b100000000;
assign racing[12][11] = 9'b100000000;
assign racing[12][12] = 9'b100000000;
assign racing[12][13] = 9'b100000000;
assign racing[12][14] = 9'b100000000;
assign racing[12][15] = 9'b100000000;
assign racing[12][16] = 9'b100000000;
assign racing[12][17] = 9'b100100100;
assign racing[12][18] = 9'b100101001;
assign racing[12][19] = 9'b100101001;
assign racing[12][20] = 9'b101001001;
assign racing[12][21] = 9'b100101001;
assign racing[13][4] = 9'b100100100;
assign racing[13][5] = 9'b101001001;
assign racing[13][6] = 9'b101001001;
assign racing[13][7] = 9'b100101001;
assign racing[13][8] = 9'b100100100;
assign racing[13][9] = 9'b100100100;
assign racing[13][10] = 9'b100100100;
assign racing[13][11] = 9'b100100100;
assign racing[13][12] = 9'b100100100;
assign racing[13][13] = 9'b100100100;
assign racing[13][14] = 9'b100100100;
assign racing[13][15] = 9'b100100100;
assign racing[13][16] = 9'b100100100;
assign racing[13][17] = 9'b100100100;
assign racing[13][18] = 9'b100101001;
assign racing[13][19] = 9'b100101001;
assign racing[13][20] = 9'b101001001;
assign racing[13][21] = 9'b100101001;
assign racing[14][4] = 9'b100100100;
assign racing[14][5] = 9'b101001001;
assign racing[14][6] = 9'b100101001;
assign racing[14][7] = 9'b100101001;
assign racing[14][8] = 9'b100101001;
assign racing[14][9] = 9'b100101001;
assign racing[14][10] = 9'b100101001;
assign racing[14][11] = 9'b100101001;
assign racing[14][12] = 9'b100101001;
assign racing[14][13] = 9'b100101001;
assign racing[14][14] = 9'b100101001;
assign racing[14][15] = 9'b100101001;
assign racing[14][16] = 9'b100101001;
assign racing[14][17] = 9'b100101001;
assign racing[14][18] = 9'b100101001;
assign racing[14][19] = 9'b100101001;
assign racing[14][20] = 9'b100101001;
assign racing[14][21] = 9'b100101001;
assign racing[15][4] = 9'b100100100;
assign racing[15][5] = 9'b100101001;
assign racing[15][6] = 9'b100101001;
assign racing[15][7] = 9'b100101001;
assign racing[15][8] = 9'b100101001;
assign racing[15][9] = 9'b100101001;
assign racing[15][10] = 9'b100101001;
assign racing[15][11] = 9'b100101001;
assign racing[15][12] = 9'b100101001;
assign racing[15][13] = 9'b100101001;
assign racing[15][14] = 9'b100101001;
assign racing[15][15] = 9'b100101001;
assign racing[15][16] = 9'b100101001;
assign racing[15][17] = 9'b100101001;
assign racing[15][18] = 9'b100101001;
assign racing[15][19] = 9'b100100101;
assign racing[15][20] = 9'b100101001;
assign racing[15][21] = 9'b100101001;
assign racing[16][4] = 9'b100100100;
assign racing[16][5] = 9'b100101001;
assign racing[16][6] = 9'b100100100;
assign racing[16][7] = 9'b100100101;
assign racing[16][8] = 9'b100101001;
assign racing[16][9] = 9'b100101001;
assign racing[16][10] = 9'b100101001;
assign racing[16][11] = 9'b100101001;
assign racing[16][12] = 9'b100101001;
assign racing[16][13] = 9'b100101001;
assign racing[16][14] = 9'b100101001;
assign racing[16][15] = 9'b100101001;
assign racing[16][16] = 9'b100101001;
assign racing[16][17] = 9'b100101001;
assign racing[16][18] = 9'b100101001;
assign racing[16][19] = 9'b100100100;
assign racing[16][20] = 9'b100101001;
assign racing[16][21] = 9'b100101001;
assign racing[17][4] = 9'b100100100;
assign racing[17][5] = 9'b100101001;
assign racing[17][6] = 9'b100100100;
assign racing[17][7] = 9'b100101001;
assign racing[17][8] = 9'b100101001;
assign racing[17][9] = 9'b100101001;
assign racing[17][10] = 9'b100101001;
assign racing[17][11] = 9'b100101001;
assign racing[17][12] = 9'b100101001;
assign racing[17][13] = 9'b100101001;
assign racing[17][14] = 9'b100101001;
assign racing[17][15] = 9'b101001001;
assign racing[17][16] = 9'b101001001;
assign racing[17][17] = 9'b100101001;
assign racing[17][18] = 9'b100101001;
assign racing[17][19] = 9'b100100100;
assign racing[17][20] = 9'b100101001;
assign racing[17][21] = 9'b100101001;
assign racing[18][4] = 9'b100000000;
assign racing[18][5] = 9'b100101001;
assign racing[18][6] = 9'b100100100;
assign racing[18][7] = 9'b100101001;
assign racing[18][8] = 9'b100101001;
assign racing[18][9] = 9'b100101001;
assign racing[18][10] = 9'b100101001;
assign racing[18][11] = 9'b100101001;
assign racing[18][12] = 9'b100101001;
assign racing[18][13] = 9'b100101001;
assign racing[18][14] = 9'b101001001;
assign racing[18][15] = 9'b101001001;
assign racing[18][16] = 9'b101001001;
assign racing[18][17] = 9'b100101001;
assign racing[18][18] = 9'b100101001;
assign racing[18][19] = 9'b100100100;
assign racing[18][20] = 9'b100100100;
assign racing[18][21] = 9'b100101001;
assign racing[19][5] = 9'b100100100;
assign racing[19][6] = 9'b100100100;
assign racing[19][7] = 9'b100101001;
assign racing[19][8] = 9'b100101001;
assign racing[19][9] = 9'b100101001;
assign racing[19][10] = 9'b100101001;
assign racing[19][11] = 9'b100101001;
assign racing[19][12] = 9'b100101001;
assign racing[19][13] = 9'b101001001;
assign racing[19][14] = 9'b101001001;
assign racing[19][15] = 9'b101001001;
assign racing[19][16] = 9'b101001001;
assign racing[19][17] = 9'b101001001;
assign racing[19][18] = 9'b100101001;
assign racing[19][19] = 9'b100100100;
assign racing[19][20] = 9'b100100100;
assign racing[19][21] = 9'b100101001;
assign racing[20][5] = 9'b100100100;
assign racing[20][6] = 9'b100100100;
assign racing[20][7] = 9'b100101001;
assign racing[20][8] = 9'b100101001;
assign racing[20][9] = 9'b100101001;
assign racing[20][10] = 9'b100101001;
assign racing[20][11] = 9'b100101001;
assign racing[20][12] = 9'b101001001;
assign racing[20][13] = 9'b101001001;
assign racing[20][14] = 9'b101001001;
assign racing[20][15] = 9'b101001001;
assign racing[20][16] = 9'b101001001;
assign racing[20][17] = 9'b101001001;
assign racing[20][18] = 9'b100101001;
assign racing[20][19] = 9'b100100100;
assign racing[20][20] = 9'b100100100;
assign racing[20][21] = 9'b100101001;
assign racing[21][5] = 9'b100100100;
assign racing[21][6] = 9'b100100100;
assign racing[21][7] = 9'b100101001;
assign racing[21][8] = 9'b100101001;
assign racing[21][9] = 9'b100101001;
assign racing[21][10] = 9'b100101001;
assign racing[21][11] = 9'b100101001;
assign racing[21][12] = 9'b101001001;
assign racing[21][13] = 9'b101001001;
assign racing[21][14] = 9'b101001001;
assign racing[21][15] = 9'b101001001;
assign racing[21][16] = 9'b101001001;
assign racing[21][17] = 9'b101001001;
assign racing[21][18] = 9'b100101001;
assign racing[21][19] = 9'b100100100;
assign racing[21][20] = 9'b100100100;
assign racing[21][21] = 9'b100101001;
assign racing[22][5] = 9'b100100100;
assign racing[22][6] = 9'b100100100;
assign racing[22][7] = 9'b100101001;
assign racing[22][8] = 9'b100101001;
assign racing[22][9] = 9'b100101001;
assign racing[22][10] = 9'b100101001;
assign racing[22][11] = 9'b101001001;
assign racing[22][12] = 9'b101001001;
assign racing[22][13] = 9'b101001001;
assign racing[22][14] = 9'b101001001;
assign racing[22][15] = 9'b101001001;
assign racing[22][16] = 9'b101001001;
assign racing[22][17] = 9'b101001001;
assign racing[22][18] = 9'b100101001;
assign racing[22][19] = 9'b100100100;
assign racing[22][20] = 9'b100100100;
assign racing[22][21] = 9'b100101001;
assign racing[23][5] = 9'b100100100;
assign racing[23][6] = 9'b100100100;
assign racing[23][7] = 9'b100101001;
assign racing[23][8] = 9'b100101001;
assign racing[23][9] = 9'b100101001;
assign racing[23][10] = 9'b100101001;
assign racing[23][11] = 9'b101001001;
assign racing[23][12] = 9'b101001001;
assign racing[23][13] = 9'b101001001;
assign racing[23][14] = 9'b101001001;
assign racing[23][15] = 9'b101001001;
assign racing[23][16] = 9'b101001001;
assign racing[23][17] = 9'b101001001;
assign racing[23][18] = 9'b100101001;
assign racing[23][19] = 9'b100100100;
assign racing[23][20] = 9'b100100100;
assign racing[23][21] = 9'b100101001;
assign racing[24][5] = 9'b100100100;
assign racing[24][6] = 9'b100100100;
assign racing[24][7] = 9'b100101001;
assign racing[24][8] = 9'b100101001;
assign racing[24][9] = 9'b100101001;
assign racing[24][10] = 9'b100101001;
assign racing[24][11] = 9'b101001001;
assign racing[24][12] = 9'b101001001;
assign racing[24][13] = 9'b101001001;
assign racing[24][14] = 9'b101001001;
assign racing[24][15] = 9'b101001001;
assign racing[24][16] = 9'b101001001;
assign racing[24][17] = 9'b101001001;
assign racing[24][18] = 9'b100101001;
assign racing[24][19] = 9'b100100100;
assign racing[24][20] = 9'b100100100;
assign racing[25][5] = 9'b100100100;
assign racing[25][6] = 9'b100100100;
assign racing[25][7] = 9'b100101001;
assign racing[25][8] = 9'b100101001;
assign racing[25][9] = 9'b100101001;
assign racing[25][10] = 9'b100101001;
assign racing[25][11] = 9'b101001001;
assign racing[25][12] = 9'b101001001;
assign racing[25][13] = 9'b101001001;
assign racing[25][14] = 9'b101001001;
assign racing[25][15] = 9'b101001001;
assign racing[25][16] = 9'b101001001;
assign racing[25][17] = 9'b100101001;
assign racing[25][18] = 9'b100101001;
assign racing[25][19] = 9'b100100100;
assign racing[25][20] = 9'b100100100;
assign racing[25][21] = 9'b100101001;
assign racing[26][5] = 9'b100100100;
assign racing[26][6] = 9'b100100100;
assign racing[26][7] = 9'b100100100;
assign racing[26][8] = 9'b100101001;
assign racing[26][9] = 9'b100101001;
assign racing[26][10] = 9'b100101001;
assign racing[26][11] = 9'b100101001;
assign racing[26][12] = 9'b100101001;
assign racing[26][13] = 9'b100101001;
assign racing[26][14] = 9'b100101001;
assign racing[26][15] = 9'b100101001;
assign racing[26][16] = 9'b100101001;
assign racing[26][17] = 9'b100101001;
assign racing[26][18] = 9'b100101001;
assign racing[26][19] = 9'b100100100;
assign racing[26][20] = 9'b100100100;
assign racing[26][21] = 9'b100101001;
assign racing[27][5] = 9'b100100100;
assign racing[27][6] = 9'b100100000;
assign racing[27][7] = 9'b100000000;
assign racing[27][8] = 9'b100100100;
assign racing[27][9] = 9'b100100100;
assign racing[27][10] = 9'b100100100;
assign racing[27][11] = 9'b100100100;
assign racing[27][12] = 9'b100100101;
assign racing[27][13] = 9'b100100101;
assign racing[27][14] = 9'b100100101;
assign racing[27][15] = 9'b100100100;
assign racing[27][16] = 9'b100100100;
assign racing[27][17] = 9'b100100100;
assign racing[27][18] = 9'b100100000;
assign racing[27][19] = 9'b100000000;
assign racing[27][20] = 9'b100100100;
assign racing[27][21] = 9'b100100100;
assign racing[28][2] = 9'b100100101;
assign racing[28][3] = 9'b100101001;
assign racing[28][4] = 9'b100100100;
assign racing[28][5] = 9'b100100100;
assign racing[28][6] = 9'b100000000;
assign racing[28][7] = 9'b100000000;
assign racing[28][8] = 9'b100000000;
assign racing[28][9] = 9'b100000000;
assign racing[28][10] = 9'b100000000;
assign racing[28][11] = 9'b100000000;
assign racing[28][12] = 9'b100000000;
assign racing[28][13] = 9'b100000000;
assign racing[28][14] = 9'b100000000;
assign racing[28][15] = 9'b100000000;
assign racing[28][16] = 9'b100000000;
assign racing[28][17] = 9'b100000000;
assign racing[28][18] = 9'b100000000;
assign racing[28][19] = 9'b100000000;
assign racing[28][20] = 9'b100100100;
assign racing[28][21] = 9'b100100101;
assign racing[28][22] = 9'b100100100;
assign racing[28][23] = 9'b100101001;
assign racing[29][2] = 9'b100100101;
assign racing[29][3] = 9'b101001001;
assign racing[29][4] = 9'b101001001;
assign racing[29][5] = 9'b100100101;
assign racing[29][6] = 9'b100000000;
assign racing[29][7] = 9'b100000000;
assign racing[29][8] = 9'b100000000;
assign racing[29][9] = 9'b100000000;
assign racing[29][10] = 9'b100000000;
assign racing[29][11] = 9'b100000000;
assign racing[29][12] = 9'b100000000;
assign racing[29][13] = 9'b100000000;
assign racing[29][14] = 9'b100000000;
assign racing[29][15] = 9'b100000000;
assign racing[29][16] = 9'b100000000;
assign racing[29][17] = 9'b100000000;
assign racing[29][18] = 9'b100000000;
assign racing[29][19] = 9'b100000000;
assign racing[29][20] = 9'b100100100;
assign racing[29][21] = 9'b100101001;
assign racing[29][22] = 9'b101001001;
assign racing[29][23] = 9'b100101001;
assign racing[30][4] = 9'b100100101;
assign racing[30][5] = 9'b100100101;
assign racing[30][6] = 9'b100000000;
assign racing[30][7] = 9'b100000000;
assign racing[30][8] = 9'b100000000;
assign racing[30][9] = 9'b100000000;
assign racing[30][10] = 9'b100000000;
assign racing[30][11] = 9'b100000000;
assign racing[30][12] = 9'b100000000;
assign racing[30][13] = 9'b100000000;
assign racing[30][14] = 9'b100000000;
assign racing[30][15] = 9'b100000000;
assign racing[30][16] = 9'b100000000;
assign racing[30][17] = 9'b100000000;
assign racing[30][18] = 9'b100000000;
assign racing[30][19] = 9'b100000000;
assign racing[30][20] = 9'b100100100;
assign racing[30][21] = 9'b100101001;
assign racing[30][22] = 9'b100101001;
assign racing[31][5] = 9'b100100101;
assign racing[31][6] = 9'b100100000;
assign racing[31][7] = 9'b100000000;
assign racing[31][8] = 9'b100000000;
assign racing[31][9] = 9'b100000000;
assign racing[31][10] = 9'b100000000;
assign racing[31][11] = 9'b100000000;
assign racing[31][12] = 9'b100000000;
assign racing[31][13] = 9'b100000000;
assign racing[31][14] = 9'b100000000;
assign racing[31][15] = 9'b100000000;
assign racing[31][16] = 9'b100000000;
assign racing[31][17] = 9'b100000000;
assign racing[31][18] = 9'b100000000;
assign racing[31][19] = 9'b100000000;
assign racing[31][20] = 9'b100100101;
assign racing[31][21] = 9'b100101001;
assign racing[32][4] = 9'b100000000;
assign racing[32][5] = 9'b100101001;
assign racing[32][6] = 9'b100100100;
assign racing[32][7] = 9'b100000000;
assign racing[32][8] = 9'b100000000;
assign racing[32][9] = 9'b100000000;
assign racing[32][10] = 9'b100000000;
assign racing[32][11] = 9'b100000000;
assign racing[32][12] = 9'b100000000;
assign racing[32][13] = 9'b100000000;
assign racing[32][14] = 9'b100000000;
assign racing[32][15] = 9'b100000000;
assign racing[32][16] = 9'b100000000;
assign racing[32][17] = 9'b100000000;
assign racing[32][18] = 9'b100000000;
assign racing[32][19] = 9'b100000000;
assign racing[32][20] = 9'b100100101;
assign racing[32][21] = 9'b100101001;
assign racing[33][4] = 9'b100000000;
assign racing[33][5] = 9'b100101001;
assign racing[33][6] = 9'b100100100;
assign racing[33][7] = 9'b100000000;
assign racing[33][8] = 9'b100000000;
assign racing[33][9] = 9'b100000000;
assign racing[33][10] = 9'b100000000;
assign racing[33][11] = 9'b100000000;
assign racing[33][12] = 9'b100000000;
assign racing[33][13] = 9'b100000000;
assign racing[33][14] = 9'b100000000;
assign racing[33][15] = 9'b100000000;
assign racing[33][16] = 9'b100000000;
assign racing[33][17] = 9'b100000000;
assign racing[33][18] = 9'b100000000;
assign racing[33][19] = 9'b100100100;
assign racing[33][20] = 9'b100101001;
assign racing[33][21] = 9'b100101001;
assign racing[34][4] = 9'b100000100;
assign racing[34][5] = 9'b100101001;
assign racing[34][6] = 9'b101001001;
assign racing[34][7] = 9'b100100100;
assign racing[34][8] = 9'b100000000;
assign racing[34][9] = 9'b100000000;
assign racing[34][10] = 9'b100000000;
assign racing[34][11] = 9'b100000000;
assign racing[34][12] = 9'b100000000;
assign racing[34][13] = 9'b100000000;
assign racing[34][14] = 9'b100000000;
assign racing[34][15] = 9'b100000000;
assign racing[34][16] = 9'b100000000;
assign racing[34][17] = 9'b100000000;
assign racing[34][18] = 9'b100100100;
assign racing[34][19] = 9'b101001001;
assign racing[34][20] = 9'b101001001;
assign racing[34][21] = 9'b100101001;
assign racing[35][4] = 9'b100000100;
assign racing[35][5] = 9'b100101001;
assign racing[35][6] = 9'b101001001;
assign racing[35][7] = 9'b101001001;
assign racing[35][8] = 9'b101001001;
assign racing[35][9] = 9'b100100100;
assign racing[35][10] = 9'b100100100;
assign racing[35][11] = 9'b100100100;
assign racing[35][12] = 9'b100100100;
assign racing[35][13] = 9'b100100100;
assign racing[35][14] = 9'b100100100;
assign racing[35][15] = 9'b100100100;
assign racing[35][16] = 9'b100100100;
assign racing[35][17] = 9'b101001001;
assign racing[35][18] = 9'b101001001;
assign racing[35][19] = 9'b101001001;
assign racing[35][20] = 9'b101001001;
assign racing[35][21] = 9'b100101001;
assign racing[36][4] = 9'b100000100;
assign racing[36][5] = 9'b100101001;
assign racing[36][6] = 9'b101001001;
assign racing[36][7] = 9'b101001001;
assign racing[36][8] = 9'b101001001;
assign racing[36][9] = 9'b101001001;
assign racing[36][10] = 9'b101001001;
assign racing[36][11] = 9'b101001001;
assign racing[36][12] = 9'b101001001;
assign racing[36][13] = 9'b101001001;
assign racing[36][14] = 9'b101001001;
assign racing[36][15] = 9'b101001001;
assign racing[36][16] = 9'b101001001;
assign racing[36][17] = 9'b101001001;
assign racing[36][18] = 9'b101001001;
assign racing[36][19] = 9'b101001001;
assign racing[36][20] = 9'b100101001;
assign racing[36][21] = 9'b100101001;
assign racing[37][4] = 9'b100100100;
assign racing[37][5] = 9'b100101001;
assign racing[37][6] = 9'b101001001;
assign racing[37][7] = 9'b101001001;
assign racing[37][8] = 9'b101001001;
assign racing[37][9] = 9'b101001001;
assign racing[37][10] = 9'b101001001;
assign racing[37][11] = 9'b101001001;
assign racing[37][12] = 9'b101001001;
assign racing[37][13] = 9'b101001001;
assign racing[37][14] = 9'b101001001;
assign racing[37][15] = 9'b101001001;
assign racing[37][16] = 9'b101001001;
assign racing[37][17] = 9'b101001001;
assign racing[37][18] = 9'b101001001;
assign racing[37][19] = 9'b101001001;
assign racing[37][20] = 9'b100101001;
assign racing[37][21] = 9'b100101001;
assign racing[38][4] = 9'b100100100;
assign racing[38][5] = 9'b100101001;
assign racing[38][6] = 9'b101001001;
assign racing[38][7] = 9'b101001001;
assign racing[38][8] = 9'b100100100;
assign racing[38][9] = 9'b101001001;
assign racing[38][10] = 9'b101001001;
assign racing[38][11] = 9'b101001001;
assign racing[38][12] = 9'b101001001;
assign racing[38][13] = 9'b101001001;
assign racing[38][14] = 9'b101001001;
assign racing[38][15] = 9'b101001001;
assign racing[38][16] = 9'b101001001;
assign racing[38][17] = 9'b100100100;
assign racing[38][18] = 9'b100100101;
assign racing[38][19] = 9'b101001001;
assign racing[38][20] = 9'b100101001;
assign racing[38][21] = 9'b100101001;
assign racing[39][4] = 9'b100000100;
assign racing[39][5] = 9'b100101001;
assign racing[39][6] = 9'b100101001;
assign racing[39][7] = 9'b101001001;
assign racing[39][8] = 9'b100000100;
assign racing[39][9] = 9'b100101001;
assign racing[39][10] = 9'b101001001;
assign racing[39][11] = 9'b101001001;
assign racing[39][12] = 9'b101001001;
assign racing[39][13] = 9'b101001001;
assign racing[39][14] = 9'b101001001;
assign racing[39][15] = 9'b101001001;
assign racing[39][16] = 9'b101001001;
assign racing[39][17] = 9'b100000100;
assign racing[39][18] = 9'b100101001;
assign racing[39][19] = 9'b101001001;
assign racing[39][20] = 9'b100101001;
assign racing[39][21] = 9'b100101001;
assign racing[40][4] = 9'b100000000;
assign racing[40][5] = 9'b100101001;
assign racing[40][6] = 9'b100101001;
assign racing[40][7] = 9'b101001001;
assign racing[40][8] = 9'b100100100;
assign racing[40][9] = 9'b100100101;
assign racing[40][10] = 9'b101001001;
assign racing[40][11] = 9'b101001001;
assign racing[40][12] = 9'b101001001;
assign racing[40][13] = 9'b101001001;
assign racing[40][14] = 9'b101001001;
assign racing[40][15] = 9'b101001001;
assign racing[40][16] = 9'b101001001;
assign racing[40][17] = 9'b100100100;
assign racing[40][18] = 9'b101001001;
assign racing[40][19] = 9'b101001001;
assign racing[40][20] = 9'b100101001;
assign racing[40][21] = 9'b100101001;
assign racing[41][5] = 9'b100101001;
assign racing[41][6] = 9'b100101001;
assign racing[41][7] = 9'b101001001;
assign racing[41][8] = 9'b100100101;
assign racing[41][9] = 9'b100100100;
assign racing[41][10] = 9'b101001001;
assign racing[41][11] = 9'b101001001;
assign racing[41][12] = 9'b101001001;
assign racing[41][13] = 9'b101001001;
assign racing[41][14] = 9'b101001001;
assign racing[41][15] = 9'b101001001;
assign racing[41][16] = 9'b100101001;
assign racing[41][17] = 9'b100100100;
assign racing[41][18] = 9'b101001001;
assign racing[41][19] = 9'b100101001;
assign racing[41][20] = 9'b100101001;
assign racing[41][21] = 9'b100101001;
assign racing[42][5] = 9'b100100101;
assign racing[42][6] = 9'b101001001;
assign racing[42][7] = 9'b100101001;
assign racing[42][8] = 9'b101001001;
assign racing[42][9] = 9'b100100101;
assign racing[42][10] = 9'b101001001;
assign racing[42][11] = 9'b101001001;
assign racing[42][12] = 9'b101001001;
assign racing[42][13] = 9'b101001001;
assign racing[42][14] = 9'b101001001;
assign racing[42][15] = 9'b101001001;
assign racing[42][16] = 9'b100101001;
assign racing[42][17] = 9'b100101001;
assign racing[42][18] = 9'b101001001;
assign racing[42][19] = 9'b100100101;
assign racing[42][20] = 9'b101001001;
assign racing[43][5] = 9'b100000000;
assign racing[43][6] = 9'b101101101;
assign racing[43][7] = 9'b101101101;
assign racing[43][8] = 9'b100101001;
assign racing[43][9] = 9'b101001001;
assign racing[43][10] = 9'b101001001;
assign racing[43][11] = 9'b101001001;
assign racing[43][12] = 9'b101001001;
assign racing[43][13] = 9'b101001001;
assign racing[43][14] = 9'b101001001;
assign racing[43][15] = 9'b101001001;
assign racing[43][16] = 9'b101001001;
assign racing[43][17] = 9'b100101001;
assign racing[43][18] = 9'b100100101;
assign racing[43][19] = 9'b101110001;
assign racing[43][20] = 9'b101101101;
assign racing[44][6] = 9'b101001001;
assign racing[44][7] = 9'b111111111;
assign racing[44][8] = 9'b101110001;
assign racing[44][9] = 9'b100100101;
assign racing[44][10] = 9'b100101001;
assign racing[44][11] = 9'b101001001;
assign racing[44][12] = 9'b101001001;
assign racing[44][13] = 9'b101001001;
assign racing[44][14] = 9'b101001001;
assign racing[44][15] = 9'b101001001;
assign racing[44][16] = 9'b100101001;
assign racing[44][17] = 9'b100100101;
assign racing[44][18] = 9'b110010010;
assign racing[44][19] = 9'b110110110;
assign racing[44][20] = 9'b100101001;
assign racing[45][7] = 9'b101001101;
assign racing[45][8] = 9'b111111111;
assign racing[45][9] = 9'b101001001;
assign racing[45][10] = 9'b100100101;
assign racing[45][11] = 9'b100101001;
assign racing[45][12] = 9'b100101001;
assign racing[45][13] = 9'b100101001;
assign racing[45][14] = 9'b100101001;
assign racing[45][15] = 9'b100101001;
assign racing[45][16] = 9'b100100101;
assign racing[45][17] = 9'b101101101;
assign racing[45][18] = 9'b111111111;
assign racing[45][19] = 9'b101001001;
assign racing[46][8] = 9'b101101101;
assign racing[46][9] = 9'b101101101;
assign racing[46][10] = 9'b100101001;
assign racing[46][11] = 9'b100101001;
assign racing[46][12] = 9'b100101001;
assign racing[46][13] = 9'b100101001;
assign racing[46][14] = 9'b100101001;
assign racing[46][15] = 9'b100101001;
assign racing[46][16] = 9'b100101001;
assign racing[46][17] = 9'b101101101;
assign racing[46][18] = 9'b101001101;
assign racing[47][9] = 9'b100101001;
assign racing[47][10] = 9'b100101001;
assign racing[47][11] = 9'b100101001;
assign racing[47][12] = 9'b100101001;
assign racing[47][13] = 9'b100101001;
assign racing[47][14] = 9'b100101001;
assign racing[47][15] = 9'b100101001;
assign racing[47][16] = 9'b100101001;
assign racing[47][17] = 9'b100101001;
assign racing[48][12] = 9'b100101001;
assign racing[48][13] = 9'b100101001;
assign racing[48][14] = 9'b100101001;
//Total de Lineas = 764
endmodule

