`timescale 1ns / 1ps
module game_over (
input enable,
input clock,
input [9:0] posx, posy,
input [9:0] hcount,
input [9:0] vcount,
output reg[2:0] red,
output reg[2:0] green,
output reg[1:0] blue,
output reg data);

always @(posedge clock)
begin
	if(enable)
	begin
		if(hcount >= posx & hcount < posx + RESOLUCION_X & vcount >= posy & vcount < posy + RESOLUCION_Y)
		begin
			if (game_over[vcount - posy][hcount - posx][8] == 1'b1)
			begin
				red   <= game_over[vcount- posy][hcount- posx][7:5];
				green <= game_over[vcount- posy][hcount- posx][4:2];
            blue 	<= game_over[vcount- posy][hcount- posx][1:0];
				data  <= 1'b1;
			end
			else
				data <= 0;
			end
		else
		data <= 0;
	end
end

parameter RESOLUCION_X = 50;
parameter RESOLUCION_Y = 25;
wire [8:0] game_over[RESOLUCION_Y - 1'b1 : 0][RESOLUCION_X - 1'b1 : 0];
assign game_over[0][24] = 9'b100000001;
assign game_over[0][25] = 9'b100000001;
assign game_over[1][23] = 9'b100000001;
assign game_over[1][24] = 9'b100000001;
assign game_over[1][25] = 9'b100000001;
assign game_over[1][26] = 9'b100000001;
assign game_over[2][22] = 9'b100000001;
assign game_over[2][23] = 9'b100000001;
assign game_over[2][24] = 9'b100000001;
assign game_over[2][25] = 9'b100000001;
assign game_over[2][26] = 9'b100000001;
assign game_over[2][27] = 9'b100000001;
assign game_over[3][21] = 9'b100000001;
assign game_over[3][22] = 9'b100000001;
assign game_over[3][23] = 9'b100000001;
assign game_over[3][24] = 9'b100000001;
assign game_over[3][25] = 9'b100000001;
assign game_over[3][26] = 9'b100000001;
assign game_over[3][27] = 9'b100000001;
assign game_over[3][28] = 9'b100000001;
assign game_over[4][0] = 9'b100000000;
assign game_over[4][1] = 9'b100000000;
assign game_over[4][2] = 9'b100000000;
assign game_over[4][3] = 9'b100000000;
assign game_over[4][4] = 9'b100000000;
assign game_over[4][5] = 9'b100000000;
assign game_over[4][6] = 9'b100000000;
assign game_over[4][7] = 9'b100000000;
assign game_over[4][8] = 9'b100000000;
assign game_over[4][9] = 9'b100000000;
assign game_over[4][10] = 9'b100000000;
assign game_over[4][11] = 9'b100000000;
assign game_over[4][12] = 9'b100000000;
assign game_over[4][13] = 9'b100000000;
assign game_over[4][14] = 9'b100000000;
assign game_over[4][15] = 9'b100000000;
assign game_over[4][16] = 9'b100000000;
assign game_over[4][17] = 9'b100000000;
assign game_over[4][18] = 9'b100000000;
assign game_over[4][19] = 9'b100000000;
assign game_over[4][20] = 9'b100000001;
assign game_over[4][21] = 9'b100000001;
assign game_over[4][22] = 9'b100000001;
assign game_over[4][23] = 9'b100000001;
assign game_over[4][24] = 9'b100000001;
assign game_over[4][25] = 9'b100000001;
assign game_over[4][26] = 9'b100000001;
assign game_over[4][27] = 9'b100000001;
assign game_over[4][28] = 9'b100000001;
assign game_over[4][29] = 9'b100000001;
assign game_over[4][30] = 9'b100000000;
assign game_over[4][31] = 9'b100000000;
assign game_over[4][32] = 9'b100000000;
assign game_over[4][33] = 9'b100000000;
assign game_over[4][34] = 9'b100000000;
assign game_over[4][35] = 9'b100000000;
assign game_over[4][36] = 9'b100000000;
assign game_over[4][37] = 9'b100000000;
assign game_over[4][38] = 9'b100000000;
assign game_over[4][39] = 9'b100000000;
assign game_over[4][40] = 9'b100000000;
assign game_over[4][41] = 9'b100000000;
assign game_over[4][42] = 9'b100000000;
assign game_over[4][43] = 9'b100000000;
assign game_over[4][44] = 9'b100000000;
assign game_over[4][45] = 9'b100000000;
assign game_over[4][46] = 9'b100000000;
assign game_over[4][47] = 9'b100000000;
assign game_over[4][48] = 9'b100000000;
assign game_over[4][49] = 9'b100000000;
assign game_over[5][0] = 9'b100000000;
assign game_over[5][1] = 9'b100000000;
assign game_over[5][2] = 9'b100000000;
assign game_over[5][3] = 9'b100000000;
assign game_over[5][4] = 9'b100000000;
assign game_over[5][5] = 9'b100000000;
assign game_over[5][6] = 9'b100000000;
assign game_over[5][7] = 9'b100000000;
assign game_over[5][8] = 9'b100000000;
assign game_over[5][9] = 9'b100000000;
assign game_over[5][10] = 9'b100000000;
assign game_over[5][11] = 9'b100000000;
assign game_over[5][12] = 9'b100000000;
assign game_over[5][13] = 9'b100000000;
assign game_over[5][14] = 9'b100000000;
assign game_over[5][15] = 9'b100000000;
assign game_over[5][16] = 9'b100000000;
assign game_over[5][17] = 9'b100000000;
assign game_over[5][18] = 9'b100000000;
assign game_over[5][19] = 9'b100000001;
assign game_over[5][20] = 9'b100000001;
assign game_over[5][21] = 9'b100000001;
assign game_over[5][22] = 9'b100000001;
assign game_over[5][23] = 9'b100000001;
assign game_over[5][24] = 9'b110000100;
assign game_over[5][25] = 9'b110000100;
assign game_over[5][26] = 9'b100000001;
assign game_over[5][27] = 9'b100000001;
assign game_over[5][28] = 9'b100000001;
assign game_over[5][29] = 9'b100000001;
assign game_over[5][30] = 9'b100000001;
assign game_over[5][31] = 9'b100000000;
assign game_over[5][32] = 9'b100000000;
assign game_over[5][33] = 9'b100000000;
assign game_over[5][34] = 9'b100000000;
assign game_over[5][35] = 9'b100000000;
assign game_over[5][36] = 9'b100000000;
assign game_over[5][37] = 9'b100000000;
assign game_over[5][38] = 9'b100000000;
assign game_over[5][39] = 9'b100000000;
assign game_over[5][40] = 9'b100000000;
assign game_over[5][41] = 9'b100000000;
assign game_over[5][42] = 9'b100000000;
assign game_over[5][43] = 9'b100000000;
assign game_over[5][44] = 9'b100000000;
assign game_over[5][45] = 9'b100000000;
assign game_over[5][46] = 9'b100000000;
assign game_over[5][47] = 9'b100000000;
assign game_over[5][48] = 9'b100000000;
assign game_over[5][49] = 9'b100000000;
assign game_over[6][0] = 9'b100000000;
assign game_over[6][1] = 9'b100000000;
assign game_over[6][2] = 9'b100000000;
assign game_over[6][3] = 9'b100000000;
assign game_over[6][4] = 9'b100000000;
assign game_over[6][5] = 9'b100000000;
assign game_over[6][6] = 9'b100000000;
assign game_over[6][7] = 9'b100000000;
assign game_over[6][8] = 9'b100000000;
assign game_over[6][9] = 9'b100000000;
assign game_over[6][10] = 9'b100000000;
assign game_over[6][11] = 9'b100000000;
assign game_over[6][12] = 9'b100000000;
assign game_over[6][13] = 9'b100000000;
assign game_over[6][14] = 9'b100000000;
assign game_over[6][15] = 9'b100000000;
assign game_over[6][16] = 9'b100000000;
assign game_over[6][17] = 9'b100000000;
assign game_over[6][18] = 9'b100000001;
assign game_over[6][19] = 9'b100000001;
assign game_over[6][20] = 9'b100000001;
assign game_over[6][21] = 9'b100000001;
assign game_over[6][22] = 9'b100100001;
assign game_over[6][23] = 9'b110100100;
assign game_over[6][24] = 9'b111100100;
assign game_over[6][25] = 9'b111100100;
assign game_over[6][26] = 9'b111100100;
assign game_over[6][27] = 9'b100100001;
assign game_over[6][28] = 9'b100000001;
assign game_over[6][29] = 9'b100000001;
assign game_over[6][30] = 9'b100000001;
assign game_over[6][31] = 9'b100000001;
assign game_over[6][32] = 9'b100000001;
assign game_over[6][33] = 9'b100000000;
assign game_over[6][34] = 9'b100000000;
assign game_over[6][35] = 9'b100000000;
assign game_over[6][36] = 9'b100000000;
assign game_over[6][37] = 9'b100000000;
assign game_over[6][38] = 9'b100000000;
assign game_over[6][39] = 9'b100000000;
assign game_over[6][40] = 9'b100000000;
assign game_over[6][41] = 9'b100000000;
assign game_over[6][42] = 9'b100000000;
assign game_over[6][43] = 9'b100000000;
assign game_over[6][44] = 9'b100000000;
assign game_over[6][45] = 9'b100000000;
assign game_over[6][46] = 9'b100000000;
assign game_over[6][47] = 9'b100000000;
assign game_over[6][48] = 9'b100000000;
assign game_over[6][49] = 9'b100000000;
assign game_over[7][0] = 9'b100000000;
assign game_over[7][1] = 9'b100000000;
assign game_over[7][2] = 9'b100000000;
assign game_over[7][3] = 9'b100000000;
assign game_over[7][4] = 9'b100000000;
assign game_over[7][5] = 9'b100000000;
assign game_over[7][6] = 9'b100000000;
assign game_over[7][7] = 9'b100000000;
assign game_over[7][8] = 9'b100000000;
assign game_over[7][9] = 9'b100000000;
assign game_over[7][10] = 9'b100000000;
assign game_over[7][11] = 9'b100000000;
assign game_over[7][12] = 9'b100000000;
assign game_over[7][13] = 9'b100000000;
assign game_over[7][14] = 9'b100000000;
assign game_over[7][15] = 9'b100000000;
assign game_over[7][16] = 9'b100000001;
assign game_over[7][17] = 9'b100000001;
assign game_over[7][18] = 9'b100000001;
assign game_over[7][19] = 9'b100000001;
assign game_over[7][20] = 9'b100000001;
assign game_over[7][21] = 9'b100100001;
assign game_over[7][22] = 9'b111100100;
assign game_over[7][23] = 9'b111100100;
assign game_over[7][24] = 9'b111100100;
assign game_over[7][25] = 9'b111100100;
assign game_over[7][26] = 9'b111100100;
assign game_over[7][27] = 9'b111100100;
assign game_over[7][28] = 9'b100100001;
assign game_over[7][29] = 9'b100000001;
assign game_over[7][30] = 9'b100000001;
assign game_over[7][31] = 9'b100000001;
assign game_over[7][32] = 9'b100000001;
assign game_over[7][33] = 9'b100000001;
assign game_over[7][34] = 9'b100000000;
assign game_over[7][35] = 9'b100000000;
assign game_over[7][36] = 9'b100000000;
assign game_over[7][37] = 9'b100000000;
assign game_over[7][38] = 9'b100000000;
assign game_over[7][39] = 9'b100000000;
assign game_over[7][40] = 9'b100000000;
assign game_over[7][41] = 9'b100000000;
assign game_over[7][42] = 9'b100000000;
assign game_over[7][43] = 9'b100000000;
assign game_over[7][44] = 9'b100000000;
assign game_over[7][45] = 9'b100000000;
assign game_over[7][46] = 9'b100000000;
assign game_over[7][47] = 9'b100000000;
assign game_over[7][48] = 9'b100000000;
assign game_over[7][49] = 9'b100000000;
assign game_over[8][0] = 9'b100000000;
assign game_over[8][1] = 9'b100000000;
assign game_over[8][2] = 9'b100000000;
assign game_over[8][3] = 9'b100000000;
assign game_over[8][4] = 9'b100000000;
assign game_over[8][5] = 9'b100000000;
assign game_over[8][6] = 9'b100000000;
assign game_over[8][7] = 9'b100000000;
assign game_over[8][8] = 9'b100000000;
assign game_over[8][9] = 9'b100000000;
assign game_over[8][10] = 9'b100000000;
assign game_over[8][11] = 9'b100000000;
assign game_over[8][12] = 9'b100000000;
assign game_over[8][13] = 9'b100000000;
assign game_over[8][14] = 9'b100000000;
assign game_over[8][15] = 9'b100000001;
assign game_over[8][16] = 9'b100000001;
assign game_over[8][17] = 9'b100000001;
assign game_over[8][18] = 9'b100000001;
assign game_over[8][19] = 9'b100000001;
assign game_over[8][20] = 9'b101000001;
assign game_over[8][21] = 9'b111100100;
assign game_over[8][22] = 9'b111100100;
assign game_over[8][23] = 9'b111100100;
assign game_over[8][24] = 9'b111100100;
assign game_over[8][25] = 9'b111100100;
assign game_over[8][26] = 9'b111100100;
assign game_over[8][27] = 9'b111100100;
assign game_over[8][28] = 9'b111100100;
assign game_over[8][29] = 9'b101000001;
assign game_over[8][30] = 9'b100000001;
assign game_over[8][31] = 9'b100000001;
assign game_over[8][32] = 9'b100000001;
assign game_over[8][33] = 9'b100000001;
assign game_over[8][34] = 9'b100000001;
assign game_over[8][35] = 9'b100000000;
assign game_over[8][36] = 9'b100000000;
assign game_over[8][37] = 9'b100000000;
assign game_over[8][38] = 9'b100000000;
assign game_over[8][39] = 9'b100000000;
assign game_over[8][40] = 9'b100000000;
assign game_over[8][41] = 9'b100000000;
assign game_over[8][42] = 9'b100000000;
assign game_over[8][43] = 9'b100000000;
assign game_over[8][44] = 9'b100000000;
assign game_over[8][45] = 9'b100000000;
assign game_over[8][46] = 9'b100000000;
assign game_over[8][47] = 9'b100000000;
assign game_over[8][48] = 9'b100000000;
assign game_over[8][49] = 9'b100000000;
assign game_over[9][0] = 9'b100000000;
assign game_over[9][1] = 9'b100000000;
assign game_over[9][2] = 9'b100000000;
assign game_over[9][3] = 9'b100000000;
assign game_over[9][4] = 9'b100000000;
assign game_over[9][5] = 9'b100000000;
assign game_over[9][6] = 9'b100000000;
assign game_over[9][7] = 9'b100000000;
assign game_over[9][8] = 9'b100000000;
assign game_over[9][9] = 9'b100000000;
assign game_over[9][10] = 9'b100000000;
assign game_over[9][11] = 9'b100000000;
assign game_over[9][12] = 9'b100000000;
assign game_over[9][13] = 9'b100000000;
assign game_over[9][14] = 9'b100000001;
assign game_over[9][15] = 9'b100000001;
assign game_over[9][16] = 9'b100000001;
assign game_over[9][17] = 9'b100000001;
assign game_over[9][18] = 9'b100000001;
assign game_over[9][19] = 9'b101100001;
assign game_over[9][20] = 9'b111100100;
assign game_over[9][21] = 9'b111100100;
assign game_over[9][22] = 9'b111100100;
assign game_over[9][23] = 9'b111100100;
assign game_over[9][24] = 9'b111100100;
assign game_over[9][25] = 9'b111100100;
assign game_over[9][26] = 9'b111100100;
assign game_over[9][27] = 9'b111100100;
assign game_over[9][28] = 9'b111100100;
assign game_over[9][29] = 9'b111100100;
assign game_over[9][30] = 9'b101100000;
assign game_over[9][31] = 9'b100000001;
assign game_over[9][32] = 9'b100000001;
assign game_over[9][33] = 9'b100000001;
assign game_over[9][34] = 9'b100000001;
assign game_over[9][35] = 9'b100000001;
assign game_over[9][36] = 9'b100000000;
assign game_over[9][37] = 9'b100000000;
assign game_over[9][38] = 9'b100000000;
assign game_over[9][39] = 9'b100000000;
assign game_over[9][40] = 9'b100000000;
assign game_over[9][41] = 9'b100000000;
assign game_over[9][42] = 9'b100000000;
assign game_over[9][43] = 9'b100000000;
assign game_over[9][44] = 9'b100000000;
assign game_over[9][45] = 9'b100000000;
assign game_over[9][46] = 9'b100000000;
assign game_over[9][47] = 9'b100000000;
assign game_over[9][48] = 9'b100000000;
assign game_over[9][49] = 9'b100000000;
assign game_over[10][0] = 9'b100000000;
assign game_over[10][1] = 9'b100000000;
assign game_over[10][2] = 9'b100000000;
assign game_over[10][3] = 9'b100000000;
assign game_over[10][4] = 9'b100000000;
assign game_over[10][5] = 9'b100000000;
assign game_over[10][6] = 9'b101101101;
assign game_over[10][7] = 9'b110010001;
assign game_over[10][8] = 9'b110010001;
assign game_over[10][9] = 9'b100000000;
assign game_over[10][10] = 9'b101101101;
assign game_over[10][11] = 9'b110010001;
assign game_over[10][12] = 9'b110010001;
assign game_over[10][13] = 9'b100100001;
assign game_over[10][14] = 9'b101101110;
assign game_over[10][15] = 9'b110010011;
assign game_over[10][16] = 9'b110001110;
assign game_over[10][17] = 9'b110010011;
assign game_over[10][18] = 9'b110110010;
assign game_over[10][19] = 9'b111101000;
assign game_over[10][20] = 9'b111101101;
assign game_over[10][21] = 9'b111110010;
assign game_over[10][22] = 9'b111110110;
assign game_over[10][23] = 9'b111101001;
assign game_over[10][24] = 9'b111100100;
assign game_over[10][25] = 9'b111100100;
assign game_over[10][26] = 9'b111100100;
assign game_over[10][27] = 9'b111100100;
assign game_over[10][28] = 9'b111101101;
assign game_over[10][29] = 9'b111110110;
assign game_over[10][30] = 9'b111110110;
assign game_over[10][31] = 9'b110000101;
assign game_over[10][32] = 9'b101101110;
assign game_over[10][33] = 9'b101000101;
assign game_over[10][34] = 9'b100100101;
assign game_over[10][35] = 9'b110001110;
assign game_over[10][36] = 9'b100100101;
assign game_over[10][37] = 9'b110010001;
assign game_over[10][38] = 9'b110010001;
assign game_over[10][39] = 9'b101101101;
assign game_over[10][40] = 9'b100000000;
assign game_over[10][41] = 9'b110010001;
assign game_over[10][42] = 9'b110010001;
assign game_over[10][43] = 9'b101101101;
assign game_over[10][44] = 9'b100000000;
assign game_over[10][45] = 9'b100000000;
assign game_over[10][46] = 9'b100000000;
assign game_over[10][47] = 9'b100000000;
assign game_over[10][48] = 9'b100000000;
assign game_over[10][49] = 9'b100000000;
assign game_over[11][0] = 9'b100000000;
assign game_over[11][1] = 9'b100000000;
assign game_over[11][2] = 9'b100000000;
assign game_over[11][3] = 9'b100000000;
assign game_over[11][4] = 9'b100000000;
assign game_over[11][5] = 9'b100000000;
assign game_over[11][6] = 9'b111111111;
assign game_over[11][7] = 9'b101101101;
assign game_over[11][8] = 9'b110010010;
assign game_over[11][9] = 9'b100000000;
assign game_over[11][10] = 9'b111111111;
assign game_over[11][11] = 9'b110001110;
assign game_over[11][12] = 9'b111111111;
assign game_over[11][13] = 9'b101000101;
assign game_over[11][14] = 9'b111111111;
assign game_over[11][15] = 9'b101101110;
assign game_over[11][16] = 9'b111111111;
assign game_over[11][17] = 9'b111110001;
assign game_over[11][18] = 9'b111111111;
assign game_over[11][19] = 9'b111101001;
assign game_over[11][20] = 9'b111111111;
assign game_over[11][21] = 9'b111110010;
assign game_over[11][22] = 9'b111101101;
assign game_over[11][23] = 9'b111100100;
assign game_over[11][24] = 9'b111100100;
assign game_over[11][25] = 9'b111100100;
assign game_over[11][26] = 9'b111100100;
assign game_over[11][27] = 9'b111100100;
assign game_over[11][28] = 9'b111111111;
assign game_over[11][29] = 9'b111110001;
assign game_over[11][30] = 9'b111111111;
assign game_over[11][31] = 9'b111101101;
assign game_over[11][32] = 9'b111110001;
assign game_over[11][33] = 9'b110010011;
assign game_over[11][34] = 9'b101101110;
assign game_over[11][35] = 9'b110110111;
assign game_over[11][36] = 9'b100100101;
assign game_over[11][37] = 9'b111111111;
assign game_over[11][38] = 9'b101101001;
assign game_over[11][39] = 9'b100100100;
assign game_over[11][40] = 9'b100100100;
assign game_over[11][41] = 9'b111111111;
assign game_over[11][42] = 9'b101101101;
assign game_over[11][43] = 9'b111111111;
assign game_over[11][44] = 9'b100000000;
assign game_over[11][45] = 9'b100000000;
assign game_over[11][46] = 9'b100000000;
assign game_over[11][47] = 9'b100000000;
assign game_over[11][48] = 9'b100000000;
assign game_over[11][49] = 9'b100000000;
assign game_over[12][0] = 9'b100000000;
assign game_over[12][1] = 9'b100000000;
assign game_over[12][2] = 9'b100000000;
assign game_over[12][3] = 9'b100000000;
assign game_over[12][4] = 9'b100000000;
assign game_over[12][5] = 9'b100000000;
assign game_over[12][6] = 9'b110110110;
assign game_over[12][7] = 9'b101001001;
assign game_over[12][8] = 9'b110110110;
assign game_over[12][9] = 9'b100000000;
assign game_over[12][10] = 9'b110110110;
assign game_over[12][11] = 9'b111110111;
assign game_over[12][12] = 9'b111111111;
assign game_over[12][13] = 9'b100100101;
assign game_over[12][14] = 9'b111110111;
assign game_over[12][15] = 9'b100100101;
assign game_over[12][16] = 9'b110110111;
assign game_over[12][17] = 9'b111101001;
assign game_over[12][18] = 9'b111110111;
assign game_over[12][19] = 9'b111101001;
assign game_over[12][20] = 9'b111110110;
assign game_over[12][21] = 9'b111111111;
assign game_over[12][22] = 9'b111101101;
assign game_over[12][23] = 9'b111100100;
assign game_over[12][24] = 9'b111100100;
assign game_over[12][25] = 9'b111100100;
assign game_over[12][26] = 9'b111100100;
assign game_over[12][27] = 9'b111100100;
assign game_over[12][28] = 9'b111111111;
assign game_over[12][29] = 9'b111101001;
assign game_over[12][30] = 9'b111110010;
assign game_over[12][31] = 9'b111101101;
assign game_over[12][32] = 9'b111101000;
assign game_over[12][33] = 9'b111111111;
assign game_over[12][34] = 9'b110110111;
assign game_over[12][35] = 9'b101001001;
assign game_over[12][36] = 9'b100100101;
assign game_over[12][37] = 9'b111111111;
assign game_over[12][38] = 9'b110010011;
assign game_over[12][39] = 9'b100100100;
assign game_over[12][40] = 9'b100000000;
assign game_over[12][41] = 9'b111111111;
assign game_over[12][42] = 9'b110110110;
assign game_over[12][43] = 9'b110110110;
assign game_over[12][44] = 9'b100000000;
assign game_over[12][45] = 9'b100000000;
assign game_over[12][46] = 9'b100000000;
assign game_over[12][47] = 9'b100000000;
assign game_over[12][48] = 9'b100000000;
assign game_over[12][49] = 9'b100000000;
assign game_over[13][0] = 9'b100000000;
assign game_over[13][1] = 9'b100000000;
assign game_over[13][2] = 9'b100000000;
assign game_over[13][3] = 9'b100000000;
assign game_over[13][4] = 9'b100000000;
assign game_over[13][5] = 9'b100000000;
assign game_over[13][6] = 9'b111111111;
assign game_over[13][7] = 9'b101101101;
assign game_over[13][8] = 9'b111111111;
assign game_over[13][9] = 9'b100100100;
assign game_over[13][10] = 9'b111111111;
assign game_over[13][11] = 9'b101001001;
assign game_over[13][12] = 9'b111111111;
assign game_over[13][13] = 9'b101000101;
assign game_over[13][14] = 9'b111111111;
assign game_over[13][15] = 9'b101000101;
assign game_over[13][16] = 9'b111111111;
assign game_over[13][17] = 9'b111101001;
assign game_over[13][18] = 9'b111111111;
assign game_over[13][19] = 9'b111101101;
assign game_over[13][20] = 9'b111111111;
assign game_over[13][21] = 9'b111110010;
assign game_over[13][22] = 9'b111101101;
assign game_over[13][23] = 9'b111100100;
assign game_over[13][24] = 9'b111100100;
assign game_over[13][25] = 9'b111100100;
assign game_over[13][26] = 9'b111100100;
assign game_over[13][27] = 9'b111100100;
assign game_over[13][28] = 9'b111111111;
assign game_over[13][29] = 9'b111110001;
assign game_over[13][30] = 9'b111111111;
assign game_over[13][31] = 9'b111101101;
assign game_over[13][32] = 9'b110100000;
assign game_over[13][33] = 9'b111111111;
assign game_over[13][34] = 9'b111111111;
assign game_over[13][35] = 9'b100000001;
assign game_over[13][36] = 9'b101000101;
assign game_over[13][37] = 9'b111111111;
assign game_over[13][38] = 9'b101101001;
assign game_over[13][39] = 9'b100100100;
assign game_over[13][40] = 9'b100100100;
assign game_over[13][41] = 9'b111111111;
assign game_over[13][42] = 9'b100100100;
assign game_over[13][43] = 9'b111111111;
assign game_over[13][44] = 9'b100000000;
assign game_over[13][45] = 9'b100000000;
assign game_over[13][46] = 9'b100000000;
assign game_over[13][47] = 9'b100000000;
assign game_over[13][48] = 9'b100000000;
assign game_over[13][49] = 9'b100000000;
assign game_over[14][0] = 9'b100000000;
assign game_over[14][1] = 9'b100000000;
assign game_over[14][2] = 9'b100000000;
assign game_over[14][3] = 9'b100000000;
assign game_over[14][4] = 9'b100000000;
assign game_over[14][5] = 9'b100000000;
assign game_over[14][6] = 9'b101101101;
assign game_over[14][7] = 9'b110010001;
assign game_over[14][8] = 9'b110010001;
assign game_over[14][9] = 9'b100000000;
assign game_over[14][10] = 9'b101101101;
assign game_over[14][11] = 9'b100000000;
assign game_over[14][12] = 9'b101101101;
assign game_over[14][13] = 9'b100100101;
assign game_over[14][14] = 9'b101101110;
assign game_over[14][15] = 9'b100100101;
assign game_over[14][16] = 9'b101101110;
assign game_over[14][17] = 9'b100100101;
assign game_over[14][18] = 9'b110001110;
assign game_over[14][19] = 9'b111101001;
assign game_over[14][20] = 9'b111101101;
assign game_over[14][21] = 9'b111110010;
assign game_over[14][22] = 9'b111110110;
assign game_over[14][23] = 9'b111101001;
assign game_over[14][24] = 9'b111100100;
assign game_over[14][25] = 9'b111100100;
assign game_over[14][26] = 9'b111100100;
assign game_over[14][27] = 9'b111100100;
assign game_over[14][28] = 9'b111101101;
assign game_over[14][29] = 9'b111110110;
assign game_over[14][30] = 9'b111110110;
assign game_over[14][31] = 9'b110000101;
assign game_over[14][32] = 9'b100000001;
assign game_over[14][33] = 9'b101001010;
assign game_over[14][34] = 9'b101101110;
assign game_over[14][35] = 9'b100000001;
assign game_over[14][36] = 9'b100100101;
assign game_over[14][37] = 9'b110010001;
assign game_over[14][38] = 9'b110010001;
assign game_over[14][39] = 9'b101101101;
assign game_over[14][40] = 9'b100000000;
assign game_over[14][41] = 9'b101101101;
assign game_over[14][42] = 9'b100000000;
assign game_over[14][43] = 9'b101101101;
assign game_over[14][44] = 9'b100000000;
assign game_over[14][45] = 9'b100000000;
assign game_over[14][46] = 9'b100000000;
assign game_over[14][47] = 9'b100000000;
assign game_over[14][48] = 9'b100000000;
assign game_over[14][49] = 9'b100000000;
assign game_over[15][0] = 9'b100000000;
assign game_over[15][1] = 9'b100000000;
assign game_over[15][2] = 9'b100000000;
assign game_over[15][3] = 9'b100000000;
assign game_over[15][4] = 9'b100000000;
assign game_over[15][5] = 9'b100000000;
assign game_over[15][6] = 9'b100000000;
assign game_over[15][7] = 9'b100000000;
assign game_over[15][8] = 9'b100000000;
assign game_over[15][9] = 9'b100000000;
assign game_over[15][10] = 9'b100000000;
assign game_over[15][11] = 9'b100000000;
assign game_over[15][12] = 9'b100000000;
assign game_over[15][13] = 9'b100000000;
assign game_over[15][14] = 9'b100000001;
assign game_over[15][15] = 9'b100000001;
assign game_over[15][16] = 9'b100000001;
assign game_over[15][17] = 9'b100000001;
assign game_over[15][18] = 9'b100000001;
assign game_over[15][19] = 9'b101100001;
assign game_over[15][20] = 9'b111100100;
assign game_over[15][21] = 9'b111100100;
assign game_over[15][22] = 9'b111100100;
assign game_over[15][23] = 9'b111100100;
assign game_over[15][24] = 9'b111100100;
assign game_over[15][25] = 9'b111100100;
assign game_over[15][26] = 9'b111100100;
assign game_over[15][27] = 9'b111100100;
assign game_over[15][28] = 9'b111100100;
assign game_over[15][29] = 9'b111100100;
assign game_over[15][30] = 9'b101100000;
assign game_over[15][31] = 9'b100000001;
assign game_over[15][32] = 9'b100000001;
assign game_over[15][33] = 9'b100000001;
assign game_over[15][34] = 9'b100000001;
assign game_over[15][35] = 9'b100000001;
assign game_over[15][36] = 9'b100000000;
assign game_over[15][37] = 9'b100000000;
assign game_over[15][38] = 9'b100000000;
assign game_over[15][39] = 9'b100000000;
assign game_over[15][40] = 9'b100000000;
assign game_over[15][41] = 9'b100000000;
assign game_over[15][42] = 9'b100000000;
assign game_over[15][43] = 9'b100000000;
assign game_over[15][44] = 9'b100000000;
assign game_over[15][45] = 9'b100000000;
assign game_over[15][46] = 9'b100000000;
assign game_over[15][47] = 9'b100000000;
assign game_over[15][48] = 9'b100000000;
assign game_over[15][49] = 9'b100000000;
assign game_over[16][0] = 9'b100000000;
assign game_over[16][1] = 9'b100000000;
assign game_over[16][2] = 9'b100000000;
assign game_over[16][3] = 9'b100000000;
assign game_over[16][4] = 9'b100000000;
assign game_over[16][5] = 9'b100000000;
assign game_over[16][6] = 9'b100000000;
assign game_over[16][7] = 9'b100000000;
assign game_over[16][8] = 9'b100000000;
assign game_over[16][9] = 9'b100000000;
assign game_over[16][10] = 9'b100000000;
assign game_over[16][11] = 9'b100000000;
assign game_over[16][12] = 9'b100000000;
assign game_over[16][13] = 9'b100000000;
assign game_over[16][14] = 9'b100000000;
assign game_over[16][15] = 9'b100000001;
assign game_over[16][16] = 9'b100000001;
assign game_over[16][17] = 9'b100000001;
assign game_over[16][18] = 9'b100000001;
assign game_over[16][19] = 9'b100000001;
assign game_over[16][20] = 9'b101000001;
assign game_over[16][21] = 9'b111100100;
assign game_over[16][22] = 9'b111100100;
assign game_over[16][23] = 9'b111100100;
assign game_over[16][24] = 9'b111100100;
assign game_over[16][25] = 9'b111100100;
assign game_over[16][26] = 9'b111100100;
assign game_over[16][27] = 9'b111100100;
assign game_over[16][28] = 9'b111100100;
assign game_over[16][29] = 9'b101000001;
assign game_over[16][30] = 9'b100000001;
assign game_over[16][31] = 9'b100000001;
assign game_over[16][32] = 9'b100000001;
assign game_over[16][33] = 9'b100000001;
assign game_over[16][34] = 9'b100000001;
assign game_over[16][35] = 9'b100000000;
assign game_over[16][36] = 9'b100000000;
assign game_over[16][37] = 9'b100000000;
assign game_over[16][38] = 9'b100000000;
assign game_over[16][39] = 9'b100000000;
assign game_over[16][40] = 9'b100000000;
assign game_over[16][41] = 9'b100000000;
assign game_over[16][42] = 9'b100000000;
assign game_over[16][43] = 9'b100000000;
assign game_over[16][44] = 9'b100000000;
assign game_over[16][45] = 9'b100000000;
assign game_over[16][46] = 9'b100000000;
assign game_over[16][47] = 9'b100000000;
assign game_over[16][48] = 9'b100000000;
assign game_over[16][49] = 9'b100000000;
assign game_over[17][0] = 9'b100000000;
assign game_over[17][1] = 9'b100000000;
assign game_over[17][2] = 9'b100000000;
assign game_over[17][3] = 9'b100000000;
assign game_over[17][4] = 9'b100000000;
assign game_over[17][5] = 9'b100000000;
assign game_over[17][6] = 9'b100000000;
assign game_over[17][7] = 9'b100000000;
assign game_over[17][8] = 9'b100000000;
assign game_over[17][9] = 9'b100000000;
assign game_over[17][10] = 9'b100000000;
assign game_over[17][11] = 9'b100000000;
assign game_over[17][12] = 9'b100000000;
assign game_over[17][13] = 9'b100000000;
assign game_over[17][14] = 9'b100000000;
assign game_over[17][15] = 9'b100000000;
assign game_over[17][16] = 9'b100000001;
assign game_over[17][17] = 9'b100000001;
assign game_over[17][18] = 9'b100000001;
assign game_over[17][19] = 9'b100000001;
assign game_over[17][20] = 9'b100000001;
assign game_over[17][21] = 9'b100100001;
assign game_over[17][22] = 9'b111100100;
assign game_over[17][23] = 9'b111100100;
assign game_over[17][24] = 9'b111100100;
assign game_over[17][25] = 9'b111100100;
assign game_over[17][26] = 9'b111100100;
assign game_over[17][27] = 9'b111100100;
assign game_over[17][28] = 9'b100100001;
assign game_over[17][29] = 9'b100000001;
assign game_over[17][30] = 9'b100000001;
assign game_over[17][31] = 9'b100000001;
assign game_over[17][32] = 9'b100000001;
assign game_over[17][33] = 9'b100000001;
assign game_over[17][34] = 9'b100000000;
assign game_over[17][35] = 9'b100000000;
assign game_over[17][36] = 9'b100000000;
assign game_over[17][37] = 9'b100000000;
assign game_over[17][38] = 9'b100000000;
assign game_over[17][39] = 9'b100000000;
assign game_over[17][40] = 9'b100000000;
assign game_over[17][41] = 9'b100000000;
assign game_over[17][42] = 9'b100000000;
assign game_over[17][43] = 9'b100000000;
assign game_over[17][44] = 9'b100000000;
assign game_over[17][45] = 9'b100000000;
assign game_over[17][46] = 9'b100000000;
assign game_over[17][47] = 9'b100000000;
assign game_over[17][48] = 9'b100000000;
assign game_over[17][49] = 9'b100000000;
assign game_over[18][0] = 9'b100000000;
assign game_over[18][1] = 9'b100000000;
assign game_over[18][2] = 9'b100000000;
assign game_over[18][3] = 9'b100000000;
assign game_over[18][4] = 9'b100000000;
assign game_over[18][5] = 9'b100000000;
assign game_over[18][6] = 9'b100000000;
assign game_over[18][7] = 9'b100000000;
assign game_over[18][8] = 9'b100000000;
assign game_over[18][9] = 9'b100000000;
assign game_over[18][10] = 9'b100000000;
assign game_over[18][11] = 9'b100000000;
assign game_over[18][12] = 9'b100000000;
assign game_over[18][13] = 9'b100000000;
assign game_over[18][14] = 9'b100000000;
assign game_over[18][15] = 9'b100000000;
assign game_over[18][16] = 9'b100000000;
assign game_over[18][17] = 9'b100000000;
assign game_over[18][18] = 9'b100000001;
assign game_over[18][19] = 9'b100000001;
assign game_over[18][20] = 9'b100000001;
assign game_over[18][21] = 9'b100000001;
assign game_over[18][22] = 9'b100100001;
assign game_over[18][23] = 9'b110100100;
assign game_over[18][24] = 9'b111100100;
assign game_over[18][25] = 9'b111100100;
assign game_over[18][26] = 9'b111100100;
assign game_over[18][27] = 9'b100100001;
assign game_over[18][28] = 9'b100000001;
assign game_over[18][29] = 9'b100000001;
assign game_over[18][30] = 9'b100000001;
assign game_over[18][31] = 9'b100000001;
assign game_over[18][32] = 9'b100000001;
assign game_over[18][33] = 9'b100000000;
assign game_over[18][34] = 9'b100000000;
assign game_over[18][35] = 9'b100000000;
assign game_over[18][36] = 9'b100000000;
assign game_over[18][37] = 9'b100000000;
assign game_over[18][38] = 9'b100000000;
assign game_over[18][39] = 9'b100000000;
assign game_over[18][40] = 9'b100000000;
assign game_over[18][41] = 9'b100000000;
assign game_over[18][42] = 9'b100000000;
assign game_over[18][43] = 9'b100000000;
assign game_over[18][44] = 9'b100000000;
assign game_over[18][45] = 9'b100000000;
assign game_over[18][46] = 9'b100000000;
assign game_over[18][47] = 9'b100000000;
assign game_over[18][48] = 9'b100000000;
assign game_over[18][49] = 9'b100000000;
assign game_over[19][0] = 9'b100000000;
assign game_over[19][1] = 9'b100000000;
assign game_over[19][2] = 9'b100000000;
assign game_over[19][3] = 9'b100000000;
assign game_over[19][4] = 9'b100000000;
assign game_over[19][5] = 9'b100000000;
assign game_over[19][6] = 9'b100000000;
assign game_over[19][7] = 9'b100000000;
assign game_over[19][8] = 9'b100000000;
assign game_over[19][9] = 9'b100000000;
assign game_over[19][10] = 9'b100000000;
assign game_over[19][11] = 9'b100000000;
assign game_over[19][12] = 9'b100000000;
assign game_over[19][13] = 9'b100000000;
assign game_over[19][14] = 9'b100000000;
assign game_over[19][15] = 9'b100000000;
assign game_over[19][16] = 9'b100000000;
assign game_over[19][17] = 9'b100000000;
assign game_over[19][18] = 9'b100000000;
assign game_over[19][19] = 9'b100000001;
assign game_over[19][20] = 9'b100000001;
assign game_over[19][21] = 9'b100000001;
assign game_over[19][22] = 9'b100000001;
assign game_over[19][23] = 9'b100000001;
assign game_over[19][24] = 9'b110000100;
assign game_over[19][25] = 9'b110000100;
assign game_over[19][26] = 9'b100000001;
assign game_over[19][27] = 9'b100000001;
assign game_over[19][28] = 9'b100000001;
assign game_over[19][29] = 9'b100000001;
assign game_over[19][30] = 9'b100000001;
assign game_over[19][31] = 9'b100000000;
assign game_over[19][32] = 9'b100000000;
assign game_over[19][33] = 9'b100000000;
assign game_over[19][34] = 9'b100000000;
assign game_over[19][35] = 9'b100000000;
assign game_over[19][36] = 9'b100000000;
assign game_over[19][37] = 9'b100000000;
assign game_over[19][38] = 9'b100000000;
assign game_over[19][39] = 9'b100000000;
assign game_over[19][40] = 9'b100000000;
assign game_over[19][41] = 9'b100000000;
assign game_over[19][42] = 9'b100000000;
assign game_over[19][43] = 9'b100000000;
assign game_over[19][44] = 9'b100000000;
assign game_over[19][45] = 9'b100000000;
assign game_over[19][46] = 9'b100000000;
assign game_over[19][47] = 9'b100000000;
assign game_over[19][48] = 9'b100000000;
assign game_over[19][49] = 9'b100000000;
assign game_over[20][0] = 9'b100000000;
assign game_over[20][1] = 9'b100000000;
assign game_over[20][2] = 9'b100000000;
assign game_over[20][3] = 9'b100000000;
assign game_over[20][4] = 9'b100000000;
assign game_over[20][5] = 9'b100000000;
assign game_over[20][6] = 9'b100000000;
assign game_over[20][7] = 9'b100000000;
assign game_over[20][8] = 9'b100000000;
assign game_over[20][9] = 9'b100000000;
assign game_over[20][10] = 9'b100000000;
assign game_over[20][11] = 9'b100000000;
assign game_over[20][12] = 9'b100000000;
assign game_over[20][13] = 9'b100000000;
assign game_over[20][14] = 9'b100000000;
assign game_over[20][15] = 9'b100000000;
assign game_over[20][16] = 9'b100000000;
assign game_over[20][17] = 9'b100000000;
assign game_over[20][18] = 9'b100000000;
assign game_over[20][19] = 9'b100000000;
assign game_over[20][20] = 9'b100000001;
assign game_over[20][21] = 9'b100000001;
assign game_over[20][22] = 9'b100000001;
assign game_over[20][23] = 9'b100000001;
assign game_over[20][24] = 9'b100000001;
assign game_over[20][25] = 9'b100000001;
assign game_over[20][26] = 9'b100000001;
assign game_over[20][27] = 9'b100000001;
assign game_over[20][28] = 9'b100000001;
assign game_over[20][29] = 9'b100000001;
assign game_over[20][30] = 9'b100000000;
assign game_over[20][31] = 9'b100000000;
assign game_over[20][32] = 9'b100000000;
assign game_over[20][33] = 9'b100000000;
assign game_over[20][34] = 9'b100000000;
assign game_over[20][35] = 9'b100000000;
assign game_over[20][36] = 9'b100000000;
assign game_over[20][37] = 9'b100000000;
assign game_over[20][38] = 9'b100000000;
assign game_over[20][39] = 9'b100000000;
assign game_over[20][40] = 9'b100000000;
assign game_over[20][41] = 9'b100000000;
assign game_over[20][42] = 9'b100000000;
assign game_over[20][43] = 9'b100000000;
assign game_over[20][44] = 9'b100000000;
assign game_over[20][45] = 9'b100000000;
assign game_over[20][46] = 9'b100000000;
assign game_over[20][47] = 9'b100000000;
assign game_over[20][48] = 9'b100000000;
assign game_over[20][49] = 9'b100000000;
assign game_over[21][21] = 9'b100000001;
assign game_over[21][22] = 9'b100000001;
assign game_over[21][23] = 9'b100000001;
assign game_over[21][24] = 9'b100000001;
assign game_over[21][25] = 9'b100000001;
assign game_over[21][26] = 9'b100000001;
assign game_over[21][27] = 9'b100000001;
assign game_over[21][28] = 9'b100000001;
assign game_over[22][22] = 9'b100000001;
assign game_over[22][23] = 9'b100000001;
assign game_over[22][24] = 9'b100000001;
assign game_over[22][25] = 9'b100000001;
assign game_over[22][26] = 9'b100000001;
assign game_over[22][27] = 9'b100000001;
assign game_over[23][23] = 9'b100000001;
assign game_over[23][24] = 9'b100000001;
assign game_over[23][25] = 9'b100000001;
assign game_over[23][26] = 9'b100000001;
assign game_over[24][24] = 9'b100000001;
assign game_over[24][25] = 9'b100000001;
//Total de Lineas = 890
endmodule

