`timescale 1ns / 1ps
module logo (
input enable,
input clock,
input [9:0] posx, posy,
input [9:0] hcount,
input [9:0] vcount,
output reg[2:0] red,
output reg[2:0] green,
output reg[1:0] blue,
output reg data);

always @(posedge clock)
begin
	if(enable)
	begin
		if(hcount >= posx & hcount < posx + RESOLUCION_X & vcount >= posy & vcount < posy + RESOLUCION_Y)
		begin
			if (logo[vcount - posy][hcount - posx][8] == 1'b1)
			begin
				red   <= logo[vcount- posy][hcount- posx][7:5];
				green <= logo[vcount- posy][hcount- posx][4:2];
            blue 	<= logo[vcount- posy][hcount- posx][1:0];
				data  <= 1'b1;
			end
			else
				data <= 0;
			end
		else
		data <= 0;
	end
end

parameter RESOLUCION_X = 100;
parameter RESOLUCION_Y = 50;
wire [8:0] logo[RESOLUCION_Y - 1'b1 : 0][RESOLUCION_X - 1'b1 : 0];
assign logo[17][35] = 9'b111111111;
assign logo[17][36] = 9'b111111111;
assign logo[17][37] = 9'b111111111;
assign logo[17][92] = 9'b111111111;
assign logo[17][93] = 9'b111111111;
assign logo[18][3] = 9'b111111111;
assign logo[18][4] = 9'b111111111;
assign logo[18][5] = 9'b111111111;
assign logo[18][6] = 9'b111111111;
assign logo[18][7] = 9'b111111111;
assign logo[18][8] = 9'b111111111;
assign logo[18][10] = 9'b111111111;
assign logo[18][11] = 9'b111111111;
assign logo[18][14] = 9'b111111111;
assign logo[18][15] = 9'b111111111;
assign logo[18][16] = 9'b111111111;
assign logo[18][18] = 9'b111111111;
assign logo[18][19] = 9'b111111111;
assign logo[18][20] = 9'b111111111;
assign logo[18][21] = 9'b111111111;
assign logo[18][22] = 9'b111111111;
assign logo[18][23] = 9'b111111111;
assign logo[18][24] = 9'b111111111;
assign logo[18][25] = 9'b111111111;
assign logo[18][28] = 9'b111111111;
assign logo[18][29] = 9'b111111111;
assign logo[18][30] = 9'b111111111;
assign logo[18][34] = 9'b111111111;
assign logo[18][35] = 9'b111111111;
assign logo[18][36] = 9'b111111111;
assign logo[18][37] = 9'b111111111;
assign logo[18][38] = 9'b111111111;
assign logo[18][41] = 9'b111111111;
assign logo[18][42] = 9'b111111111;
assign logo[18][43] = 9'b111111111;
assign logo[18][45] = 9'b111111111;
assign logo[18][46] = 9'b111111111;
assign logo[18][47] = 9'b111111111;
assign logo[18][53] = 9'b111111111;
assign logo[18][54] = 9'b111111111;
assign logo[18][55] = 9'b111111111;
assign logo[18][57] = 9'b111111111;
assign logo[18][58] = 9'b111111111;
assign logo[18][59] = 9'b111111111;
assign logo[18][61] = 9'b111111111;
assign logo[18][62] = 9'b111111111;
assign logo[18][63] = 9'b111111111;
assign logo[18][64] = 9'b111111111;
assign logo[18][65] = 9'b111111111;
assign logo[18][68] = 9'b111111111;
assign logo[18][69] = 9'b111111111;
assign logo[18][71] = 9'b111111111;
assign logo[18][72] = 9'b111111111;
assign logo[18][73] = 9'b111111111;
assign logo[18][74] = 9'b111111111;
assign logo[18][75] = 9'b111111111;
assign logo[18][76] = 9'b111111111;
assign logo[18][78] = 9'b111111111;
assign logo[18][79] = 9'b111111111;
assign logo[18][80] = 9'b111111111;
assign logo[18][81] = 9'b111111111;
assign logo[18][82] = 9'b111111111;
assign logo[18][83] = 9'b111111111;
assign logo[18][84] = 9'b111111111;
assign logo[18][85] = 9'b111111111;
assign logo[18][91] = 9'b111111111;
assign logo[18][92] = 9'b111111111;
assign logo[18][93] = 9'b111111111;
assign logo[18][94] = 9'b111111111;
assign logo[18][95] = 9'b111111111;
assign logo[19][3] = 9'b111111111;
assign logo[19][4] = 9'b111111111;
assign logo[19][5] = 9'b111111111;
assign logo[19][6] = 9'b111111111;
assign logo[19][7] = 9'b111111111;
assign logo[19][8] = 9'b111111111;
assign logo[19][10] = 9'b111111111;
assign logo[19][11] = 9'b111111111;
assign logo[19][14] = 9'b111111111;
assign logo[19][15] = 9'b111111111;
assign logo[19][16] = 9'b111111111;
assign logo[19][18] = 9'b111111111;
assign logo[19][19] = 9'b111111111;
assign logo[19][20] = 9'b111111111;
assign logo[19][21] = 9'b111111111;
assign logo[19][22] = 9'b111111111;
assign logo[19][23] = 9'b111111111;
assign logo[19][24] = 9'b111111111;
assign logo[19][25] = 9'b111111111;
assign logo[19][26] = 9'b111111111;
assign logo[19][28] = 9'b111111111;
assign logo[19][29] = 9'b111111111;
assign logo[19][33] = 9'b111111111;
assign logo[19][34] = 9'b111111111;
assign logo[19][35] = 9'b111111111;
assign logo[19][36] = 9'b111111111;
assign logo[19][37] = 9'b111111111;
assign logo[19][38] = 9'b111111111;
assign logo[19][39] = 9'b111111111;
assign logo[19][41] = 9'b111111111;
assign logo[19][42] = 9'b111111111;
assign logo[19][43] = 9'b111111111;
assign logo[19][45] = 9'b111111111;
assign logo[19][46] = 9'b111111111;
assign logo[19][47] = 9'b111111111;
assign logo[19][53] = 9'b111111111;
assign logo[19][54] = 9'b111111111;
assign logo[19][55] = 9'b111111111;
assign logo[19][57] = 9'b111111111;
assign logo[19][58] = 9'b111111111;
assign logo[19][59] = 9'b111111111;
assign logo[19][61] = 9'b111111111;
assign logo[19][62] = 9'b111111111;
assign logo[19][63] = 9'b111111111;
assign logo[19][64] = 9'b111111111;
assign logo[19][65] = 9'b111111111;
assign logo[19][68] = 9'b111111111;
assign logo[19][69] = 9'b111111111;
assign logo[19][71] = 9'b111111111;
assign logo[19][72] = 9'b111111111;
assign logo[19][73] = 9'b111111111;
assign logo[19][74] = 9'b111111111;
assign logo[19][75] = 9'b111111111;
assign logo[19][76] = 9'b111111111;
assign logo[19][78] = 9'b111111111;
assign logo[19][79] = 9'b111111111;
assign logo[19][80] = 9'b111111111;
assign logo[19][81] = 9'b111111111;
assign logo[19][82] = 9'b111111111;
assign logo[19][83] = 9'b111111111;
assign logo[19][84] = 9'b111111111;
assign logo[19][85] = 9'b111111111;
assign logo[19][90] = 9'b111111111;
assign logo[19][91] = 9'b111111111;
assign logo[19][92] = 9'b111111111;
assign logo[19][93] = 9'b111111111;
assign logo[19][94] = 9'b111111111;
assign logo[19][95] = 9'b111111111;
assign logo[20][3] = 9'b111111111;
assign logo[20][4] = 9'b111111111;
assign logo[20][5] = 9'b111111111;
assign logo[20][10] = 9'b111111111;
assign logo[20][11] = 9'b111111111;
assign logo[20][14] = 9'b111111111;
assign logo[20][15] = 9'b111111111;
assign logo[20][16] = 9'b111111111;
assign logo[20][18] = 9'b111111111;
assign logo[20][19] = 9'b111111111;
assign logo[20][21] = 9'b111111111;
assign logo[20][22] = 9'b111111111;
assign logo[20][23] = 9'b111111111;
assign logo[20][25] = 9'b111111111;
assign logo[20][26] = 9'b111111111;
assign logo[20][27] = 9'b111111111;
assign logo[20][28] = 9'b111111111;
assign logo[20][29] = 9'b111111111;
assign logo[20][33] = 9'b111111111;
assign logo[20][34] = 9'b111111111;
assign logo[20][35] = 9'b111111111;
assign logo[20][37] = 9'b111111111;
assign logo[20][38] = 9'b111111111;
assign logo[20][39] = 9'b111111111;
assign logo[20][41] = 9'b111111111;
assign logo[20][42] = 9'b111111111;
assign logo[20][43] = 9'b111111111;
assign logo[20][44] = 9'b111111111;
assign logo[20][45] = 9'b111111111;
assign logo[20][46] = 9'b111111111;
assign logo[20][47] = 9'b111111111;
assign logo[20][53] = 9'b111111111;
assign logo[20][54] = 9'b111111111;
assign logo[20][55] = 9'b111111111;
assign logo[20][57] = 9'b111111111;
assign logo[20][58] = 9'b111111111;
assign logo[20][59] = 9'b111111111;
assign logo[20][61] = 9'b111111111;
assign logo[20][62] = 9'b111111111;
assign logo[20][63] = 9'b111111111;
assign logo[20][64] = 9'b111111111;
assign logo[20][65] = 9'b111111111;
assign logo[20][68] = 9'b111111111;
assign logo[20][69] = 9'b111111111;
assign logo[20][71] = 9'b111111111;
assign logo[20][72] = 9'b111111111;
assign logo[20][73] = 9'b111111111;
assign logo[20][78] = 9'b111111111;
assign logo[20][79] = 9'b111111111;
assign logo[20][84] = 9'b111111111;
assign logo[20][85] = 9'b111111111;
assign logo[20][90] = 9'b111111111;
assign logo[20][91] = 9'b111111111;
assign logo[20][92] = 9'b111111111;
assign logo[21][3] = 9'b111111111;
assign logo[21][4] = 9'b111111111;
assign logo[21][5] = 9'b111111111;
assign logo[21][6] = 9'b111111111;
assign logo[21][7] = 9'b111111111;
assign logo[21][10] = 9'b111111111;
assign logo[21][11] = 9'b111111111;
assign logo[21][14] = 9'b111111111;
assign logo[21][15] = 9'b111111111;
assign logo[21][16] = 9'b111111111;
assign logo[21][18] = 9'b111111111;
assign logo[21][19] = 9'b111111111;
assign logo[21][20] = 9'b111111111;
assign logo[21][21] = 9'b111111111;
assign logo[21][22] = 9'b111111111;
assign logo[21][23] = 9'b111111111;
assign logo[21][25] = 9'b111111111;
assign logo[21][26] = 9'b111111111;
assign logo[21][27] = 9'b111111111;
assign logo[21][28] = 9'b111111111;
assign logo[21][32] = 9'b111111111;
assign logo[21][33] = 9'b111111111;
assign logo[21][34] = 9'b111111111;
assign logo[21][38] = 9'b111111111;
assign logo[21][39] = 9'b111111111;
assign logo[21][40] = 9'b111111111;
assign logo[21][41] = 9'b111111111;
assign logo[21][42] = 9'b111111111;
assign logo[21][43] = 9'b111111111;
assign logo[21][44] = 9'b111111111;
assign logo[21][45] = 9'b111111111;
assign logo[21][46] = 9'b111111111;
assign logo[21][47] = 9'b111111111;
assign logo[21][54] = 9'b111111111;
assign logo[21][55] = 9'b111111111;
assign logo[21][56] = 9'b111111111;
assign logo[21][57] = 9'b111111111;
assign logo[21][58] = 9'b111111111;
assign logo[21][59] = 9'b111111111;
assign logo[21][60] = 9'b111111111;
assign logo[21][61] = 9'b111111111;
assign logo[21][62] = 9'b111111111;
assign logo[21][63] = 9'b111111111;
assign logo[21][64] = 9'b111111111;
assign logo[21][65] = 9'b111111111;
assign logo[21][66] = 9'b111111111;
assign logo[21][67] = 9'b111111111;
assign logo[21][68] = 9'b111111111;
assign logo[21][69] = 9'b111111111;
assign logo[21][71] = 9'b111111111;
assign logo[21][72] = 9'b111111111;
assign logo[21][73] = 9'b111111111;
assign logo[21][74] = 9'b111111111;
assign logo[21][75] = 9'b111111111;
assign logo[21][76] = 9'b111111111;
assign logo[21][78] = 9'b111111111;
assign logo[21][79] = 9'b111111111;
assign logo[21][80] = 9'b111111111;
assign logo[21][81] = 9'b111111111;
assign logo[21][82] = 9'b111111111;
assign logo[21][84] = 9'b111111111;
assign logo[21][85] = 9'b111111111;
assign logo[21][90] = 9'b111111111;
assign logo[21][91] = 9'b111111111;
assign logo[21][92] = 9'b111111111;
assign logo[21][93] = 9'b111111111;
assign logo[21][94] = 9'b111111111;
assign logo[22][3] = 9'b111111111;
assign logo[22][4] = 9'b111111111;
assign logo[22][5] = 9'b111111111;
assign logo[22][6] = 9'b111111111;
assign logo[22][7] = 9'b111111111;
assign logo[22][8] = 9'b111111111;
assign logo[22][10] = 9'b111111111;
assign logo[22][11] = 9'b111111111;
assign logo[22][14] = 9'b111111111;
assign logo[22][15] = 9'b111111111;
assign logo[22][16] = 9'b111111111;
assign logo[22][18] = 9'b111111111;
assign logo[22][19] = 9'b111111111;
assign logo[22][20] = 9'b111111111;
assign logo[22][21] = 9'b111111111;
assign logo[22][22] = 9'b111111111;
assign logo[22][23] = 9'b111111111;
assign logo[22][26] = 9'b111111111;
assign logo[22][27] = 9'b111111111;
assign logo[22][28] = 9'b111111111;
assign logo[22][32] = 9'b111111111;
assign logo[22][33] = 9'b111111111;
assign logo[22][34] = 9'b111111111;
assign logo[22][38] = 9'b111111111;
assign logo[22][39] = 9'b111111111;
assign logo[22][40] = 9'b111111111;
assign logo[22][41] = 9'b111111111;
assign logo[22][42] = 9'b111111111;
assign logo[22][43] = 9'b111111111;
assign logo[22][44] = 9'b111111111;
assign logo[22][45] = 9'b111111111;
assign logo[22][46] = 9'b111111111;
assign logo[22][47] = 9'b111111111;
assign logo[22][54] = 9'b111111111;
assign logo[22][55] = 9'b111111111;
assign logo[22][56] = 9'b111111111;
assign logo[22][57] = 9'b111111111;
assign logo[22][58] = 9'b111111111;
assign logo[22][59] = 9'b111111111;
assign logo[22][60] = 9'b111111111;
assign logo[22][61] = 9'b111111111;
assign logo[22][62] = 9'b111111111;
assign logo[22][63] = 9'b111111111;
assign logo[22][64] = 9'b111111111;
assign logo[22][65] = 9'b111111111;
assign logo[22][66] = 9'b111111111;
assign logo[22][67] = 9'b111111111;
assign logo[22][68] = 9'b111111111;
assign logo[22][69] = 9'b111111111;
assign logo[22][71] = 9'b111111111;
assign logo[22][72] = 9'b111111111;
assign logo[22][73] = 9'b111111111;
assign logo[22][74] = 9'b111111111;
assign logo[22][75] = 9'b111111111;
assign logo[22][76] = 9'b111111111;
assign logo[22][78] = 9'b111111111;
assign logo[22][79] = 9'b111111111;
assign logo[22][80] = 9'b111111111;
assign logo[22][81] = 9'b111111111;
assign logo[22][82] = 9'b111111111;
assign logo[22][84] = 9'b111111111;
assign logo[22][85] = 9'b111111111;
assign logo[22][91] = 9'b111111111;
assign logo[22][92] = 9'b111111111;
assign logo[22][93] = 9'b111111111;
assign logo[22][94] = 9'b111111111;
assign logo[22][95] = 9'b111111111;
assign logo[23][3] = 9'b111111111;
assign logo[23][4] = 9'b111111111;
assign logo[23][5] = 9'b111111111;
assign logo[23][6] = 9'b111111111;
assign logo[23][7] = 9'b111111111;
assign logo[23][8] = 9'b111111111;
assign logo[23][10] = 9'b111111111;
assign logo[23][11] = 9'b111111111;
assign logo[23][14] = 9'b111111111;
assign logo[23][15] = 9'b111111111;
assign logo[23][16] = 9'b111111111;
assign logo[23][18] = 9'b111111111;
assign logo[23][19] = 9'b111111111;
assign logo[23][20] = 9'b111111111;
assign logo[23][21] = 9'b111111111;
assign logo[23][22] = 9'b111111111;
assign logo[23][26] = 9'b111111111;
assign logo[23][27] = 9'b111111111;
assign logo[23][32] = 9'b111111111;
assign logo[23][33] = 9'b111111111;
assign logo[23][34] = 9'b111111111;
assign logo[23][38] = 9'b111111111;
assign logo[23][39] = 9'b111111111;
assign logo[23][40] = 9'b111111111;
assign logo[23][41] = 9'b111111111;
assign logo[23][42] = 9'b111111111;
assign logo[23][43] = 9'b111111111;
assign logo[23][44] = 9'b111111111;
assign logo[23][45] = 9'b111111111;
assign logo[23][46] = 9'b111111111;
assign logo[23][47] = 9'b111111111;
assign logo[23][54] = 9'b111111111;
assign logo[23][55] = 9'b111111111;
assign logo[23][56] = 9'b111111111;
assign logo[23][57] = 9'b111111111;
assign logo[23][58] = 9'b111111111;
assign logo[23][59] = 9'b111111111;
assign logo[23][60] = 9'b111111111;
assign logo[23][61] = 9'b111111111;
assign logo[23][62] = 9'b111111111;
assign logo[23][63] = 9'b111111111;
assign logo[23][64] = 9'b111111111;
assign logo[23][65] = 9'b111111111;
assign logo[23][66] = 9'b111111111;
assign logo[23][67] = 9'b111111111;
assign logo[23][68] = 9'b111111111;
assign logo[23][69] = 9'b111111111;
assign logo[23][71] = 9'b111111111;
assign logo[23][72] = 9'b111111111;
assign logo[23][73] = 9'b111111111;
assign logo[23][74] = 9'b111111111;
assign logo[23][75] = 9'b111111111;
assign logo[23][78] = 9'b111111111;
assign logo[23][79] = 9'b111111111;
assign logo[23][80] = 9'b111111111;
assign logo[23][81] = 9'b111111111;
assign logo[23][82] = 9'b111111111;
assign logo[23][84] = 9'b111111111;
assign logo[23][85] = 9'b111111111;
assign logo[23][94] = 9'b111111111;
assign logo[23][95] = 9'b111111111;
assign logo[23][96] = 9'b111111111;
assign logo[24][3] = 9'b111111111;
assign logo[24][4] = 9'b111111111;
assign logo[24][5] = 9'b111111111;
assign logo[24][10] = 9'b111111111;
assign logo[24][11] = 9'b111111111;
assign logo[24][12] = 9'b111111111;
assign logo[24][13] = 9'b111111111;
assign logo[24][14] = 9'b111111111;
assign logo[24][15] = 9'b111111111;
assign logo[24][16] = 9'b111111111;
assign logo[24][18] = 9'b111111111;
assign logo[24][19] = 9'b111111111;
assign logo[24][21] = 9'b111111111;
assign logo[24][22] = 9'b111111111;
assign logo[24][26] = 9'b111111111;
assign logo[24][27] = 9'b111111111;
assign logo[24][33] = 9'b111111111;
assign logo[24][34] = 9'b111111111;
assign logo[24][35] = 9'b111111111;
assign logo[24][36] = 9'b111111111;
assign logo[24][37] = 9'b111111111;
assign logo[24][38] = 9'b111111111;
assign logo[24][39] = 9'b111111111;
assign logo[24][41] = 9'b111111111;
assign logo[24][42] = 9'b111111111;
assign logo[24][43] = 9'b111111111;
assign logo[24][44] = 9'b111111111;
assign logo[24][45] = 9'b111111111;
assign logo[24][46] = 9'b111111111;
assign logo[24][47] = 9'b111111111;
assign logo[24][54] = 9'b111111111;
assign logo[24][55] = 9'b111111111;
assign logo[24][56] = 9'b111111111;
assign logo[24][57] = 9'b111111111;
assign logo[24][58] = 9'b111111111;
assign logo[24][59] = 9'b111111111;
assign logo[24][60] = 9'b111111111;
assign logo[24][61] = 9'b111111111;
assign logo[24][63] = 9'b111111111;
assign logo[24][64] = 9'b111111111;
assign logo[24][65] = 9'b111111111;
assign logo[24][68] = 9'b111111111;
assign logo[24][69] = 9'b111111111;
assign logo[24][71] = 9'b111111111;
assign logo[24][72] = 9'b111111111;
assign logo[24][73] = 9'b111111111;
assign logo[24][78] = 9'b111111111;
assign logo[24][79] = 9'b111111111;
assign logo[24][80] = 9'b111111111;
assign logo[24][84] = 9'b111111111;
assign logo[24][85] = 9'b111111111;
assign logo[24][86] = 9'b111111111;
assign logo[24][87] = 9'b111111111;
assign logo[24][88] = 9'b111111111;
assign logo[24][90] = 9'b111111111;
assign logo[24][91] = 9'b111111111;
assign logo[24][92] = 9'b111111111;
assign logo[24][93] = 9'b111111111;
assign logo[24][94] = 9'b111111111;
assign logo[24][95] = 9'b111111111;
assign logo[24][96] = 9'b111111111;
assign logo[25][3] = 9'b111111111;
assign logo[25][4] = 9'b111111111;
assign logo[25][5] = 9'b111111111;
assign logo[25][10] = 9'b111111111;
assign logo[25][11] = 9'b111111111;
assign logo[25][12] = 9'b111111111;
assign logo[25][13] = 9'b111111111;
assign logo[25][14] = 9'b111111111;
assign logo[25][15] = 9'b111111111;
assign logo[25][18] = 9'b111111111;
assign logo[25][19] = 9'b111111111;
assign logo[25][21] = 9'b111111111;
assign logo[25][22] = 9'b111111111;
assign logo[25][23] = 9'b111111111;
assign logo[25][26] = 9'b111111111;
assign logo[25][27] = 9'b111111111;
assign logo[25][33] = 9'b111111111;
assign logo[25][34] = 9'b111111111;
assign logo[25][35] = 9'b111111111;
assign logo[25][36] = 9'b111111111;
assign logo[25][37] = 9'b111111111;
assign logo[25][38] = 9'b111111111;
assign logo[25][39] = 9'b111111111;
assign logo[25][41] = 9'b111111111;
assign logo[25][42] = 9'b111111111;
assign logo[25][43] = 9'b111111111;
assign logo[25][45] = 9'b111111111;
assign logo[25][46] = 9'b111111111;
assign logo[25][47] = 9'b111111111;
assign logo[25][54] = 9'b111111111;
assign logo[25][55] = 9'b111111111;
assign logo[25][56] = 9'b111111111;
assign logo[25][57] = 9'b111111111;
assign logo[25][59] = 9'b111111111;
assign logo[25][60] = 9'b111111111;
assign logo[25][61] = 9'b111111111;
assign logo[25][63] = 9'b111111111;
assign logo[25][64] = 9'b111111111;
assign logo[25][65] = 9'b111111111;
assign logo[25][68] = 9'b111111111;
assign logo[25][69] = 9'b111111111;
assign logo[25][71] = 9'b111111111;
assign logo[25][72] = 9'b111111111;
assign logo[25][73] = 9'b111111111;
assign logo[25][74] = 9'b111111111;
assign logo[25][75] = 9'b111111111;
assign logo[25][76] = 9'b111111111;
assign logo[25][78] = 9'b111111111;
assign logo[25][79] = 9'b111111111;
assign logo[25][80] = 9'b111111111;
assign logo[25][81] = 9'b111111111;
assign logo[25][82] = 9'b111111111;
assign logo[25][83] = 9'b111111111;
assign logo[25][84] = 9'b111111111;
assign logo[25][85] = 9'b111111111;
assign logo[25][86] = 9'b111111111;
assign logo[25][87] = 9'b111111111;
assign logo[25][88] = 9'b111111111;
assign logo[25][89] = 9'b111111111;
assign logo[25][90] = 9'b111111111;
assign logo[25][91] = 9'b111111111;
assign logo[25][92] = 9'b111111111;
assign logo[25][93] = 9'b111111111;
assign logo[25][94] = 9'b111111111;
assign logo[25][95] = 9'b111111111;
assign logo[26][3] = 9'b111111111;
assign logo[26][4] = 9'b111111111;
assign logo[26][5] = 9'b111111111;
assign logo[26][11] = 9'b111111111;
assign logo[26][12] = 9'b111111111;
assign logo[26][13] = 9'b111111111;
assign logo[26][14] = 9'b111111111;
assign logo[26][18] = 9'b111111111;
assign logo[26][19] = 9'b111111111;
assign logo[26][22] = 9'b111111111;
assign logo[26][23] = 9'b111111111;
assign logo[26][26] = 9'b111111111;
assign logo[26][27] = 9'b111111111;
assign logo[26][35] = 9'b111111111;
assign logo[26][36] = 9'b111111111;
assign logo[26][37] = 9'b111111111;
assign logo[26][41] = 9'b111111111;
assign logo[26][42] = 9'b111111111;
assign logo[26][43] = 9'b111111111;
assign logo[26][45] = 9'b111111111;
assign logo[26][46] = 9'b111111111;
assign logo[26][47] = 9'b111111111;
assign logo[26][55] = 9'b111111111;
assign logo[26][56] = 9'b111111111;
assign logo[26][57] = 9'b111111111;
assign logo[26][59] = 9'b111111111;
assign logo[26][60] = 9'b111111111;
assign logo[26][61] = 9'b111111111;
assign logo[26][63] = 9'b111111111;
assign logo[26][64] = 9'b111111111;
assign logo[26][65] = 9'b111111111;
assign logo[26][68] = 9'b111111111;
assign logo[26][69] = 9'b111111111;
assign logo[26][71] = 9'b111111111;
assign logo[26][72] = 9'b111111111;
assign logo[26][73] = 9'b111111111;
assign logo[26][74] = 9'b111111111;
assign logo[26][75] = 9'b111111111;
assign logo[26][76] = 9'b111111111;
assign logo[26][78] = 9'b111111111;
assign logo[26][79] = 9'b111111111;
assign logo[26][80] = 9'b111111111;
assign logo[26][81] = 9'b111111111;
assign logo[26][82] = 9'b111111111;
assign logo[26][83] = 9'b111111111;
assign logo[26][84] = 9'b111111111;
assign logo[26][85] = 9'b111111111;
assign logo[26][86] = 9'b111111111;
assign logo[26][87] = 9'b111111111;
assign logo[26][88] = 9'b111111111;
assign logo[26][89] = 9'b111111111;
assign logo[26][91] = 9'b111111111;
assign logo[26][92] = 9'b111111111;
assign logo[26][93] = 9'b111111111;
assign logo[26][94] = 9'b111111111;
//Total de Lineas = 569
endmodule

