`timescale 1ns / 1ps
module supra (
input enable,
input clock,
input [9:0] posx, posy,
input [9:0] hcount,
input [9:0] vcount,
output reg[2:0] red,
output reg[2:0] green,
output reg[1:0] blue,
output reg data);

always @(posedge clock)
begin
	if(enable)
	begin
		if(hcount >= posx & hcount < posx + RESOLUCION_X & vcount >= posy & vcount < posy + RESOLUCION_Y)
		begin
			if (supra[vcount - posy][hcount - posx][8] == 1'b1)
			begin
				red   <= supra[vcount- posy][hcount- posx][7:5];
				green <= supra[vcount- posy][hcount- posx][4:2];
            blue 	<= supra[vcount- posy][hcount- posx][1:0];
				data  <= 1'b1;
			end
			else
				data <= 0;
			end
		else
		data <= 0;
	end
end

parameter RESOLUCION_X = 20;
parameter RESOLUCION_Y = 50;
wire [8:0] supra[RESOLUCION_Y - 1'b1 : 0][RESOLUCION_X - 1'b1 : 0];
assign supra[0][4] = 9'b110000000;
assign supra[0][5] = 9'b110000000;
assign supra[0][6] = 9'b110000000;
assign supra[0][7] = 9'b110000000;
assign supra[0][8] = 9'b110000000;
assign supra[0][9] = 9'b110000000;
assign supra[0][10] = 9'b110000000;
assign supra[0][11] = 9'b110000000;
assign supra[0][12] = 9'b110000000;
assign supra[0][13] = 9'b110000000;
assign supra[0][14] = 9'b110000000;
assign supra[0][15] = 9'b110000000;
assign supra[1][3] = 9'b110000000;
assign supra[1][4] = 9'b110000100;
assign supra[1][5] = 9'b110001101;
assign supra[1][6] = 9'b110001101;
assign supra[1][7] = 9'b110100000;
assign supra[1][8] = 9'b110100000;
assign supra[1][9] = 9'b110000000;
assign supra[1][10] = 9'b110000000;
assign supra[1][11] = 9'b110100000;
assign supra[1][12] = 9'b110100000;
assign supra[1][13] = 9'b110001001;
assign supra[1][14] = 9'b110001101;
assign supra[1][15] = 9'b110000100;
assign supra[1][16] = 9'b110000000;
assign supra[2][2] = 9'b110000000;
assign supra[2][3] = 9'b110000100;
assign supra[2][4] = 9'b101111111;
assign supra[2][5] = 9'b101111111;
assign supra[2][6] = 9'b110001101;
assign supra[2][7] = 9'b110000000;
assign supra[2][8] = 9'b110000000;
assign supra[2][9] = 9'b110000000;
assign supra[2][10] = 9'b110000000;
assign supra[2][11] = 9'b110000000;
assign supra[2][12] = 9'b110000000;
assign supra[2][13] = 9'b110001101;
assign supra[2][14] = 9'b101111111;
assign supra[2][15] = 9'b101111111;
assign supra[2][16] = 9'b110000100;
assign supra[2][17] = 9'b110000000;
assign supra[3][2] = 9'b110000000;
assign supra[3][3] = 9'b110011111;
assign supra[3][4] = 9'b101111111;
assign supra[3][5] = 9'b110001101;
assign supra[3][6] = 9'b110000000;
assign supra[3][7] = 9'b110100000;
assign supra[3][8] = 9'b110100000;
assign supra[3][9] = 9'b110100000;
assign supra[3][10] = 9'b110100000;
assign supra[3][11] = 9'b110100000;
assign supra[3][12] = 9'b110100000;
assign supra[3][13] = 9'b110000000;
assign supra[3][14] = 9'b110001101;
assign supra[3][15] = 9'b101111111;
assign supra[3][16] = 9'b110011111;
assign supra[3][17] = 9'b110000100;
assign supra[4][1] = 9'b110000000;
assign supra[4][2] = 9'b110100000;
assign supra[4][3] = 9'b110001001;
assign supra[4][4] = 9'b110000000;
assign supra[4][5] = 9'b110000000;
assign supra[4][6] = 9'b110000000;
assign supra[4][7] = 9'b110100000;
assign supra[4][8] = 9'b110100000;
assign supra[4][9] = 9'b110100000;
assign supra[4][10] = 9'b110100000;
assign supra[4][11] = 9'b110100000;
assign supra[4][12] = 9'b110100000;
assign supra[4][13] = 9'b110000000;
assign supra[4][14] = 9'b110000000;
assign supra[4][15] = 9'b110000000;
assign supra[4][16] = 9'b110001001;
assign supra[4][17] = 9'b110100100;
assign supra[4][18] = 9'b110000000;
assign supra[5][1] = 9'b110000000;
assign supra[5][2] = 9'b110100000;
assign supra[5][3] = 9'b110100000;
assign supra[5][4] = 9'b110100000;
assign supra[5][5] = 9'b110000000;
assign supra[5][6] = 9'b110000000;
assign supra[5][7] = 9'b110100000;
assign supra[5][8] = 9'b110100000;
assign supra[5][9] = 9'b110100000;
assign supra[5][10] = 9'b110100000;
assign supra[5][11] = 9'b110100000;
assign supra[5][12] = 9'b110100000;
assign supra[5][13] = 9'b110000000;
assign supra[5][14] = 9'b110000000;
assign supra[5][15] = 9'b110100000;
assign supra[5][16] = 9'b110100000;
assign supra[5][17] = 9'b110100000;
assign supra[5][18] = 9'b110000000;
assign supra[6][1] = 9'b110000000;
assign supra[6][2] = 9'b110100000;
assign supra[6][3] = 9'b110000000;
assign supra[6][4] = 9'b110100000;
assign supra[6][5] = 9'b110000000;
assign supra[6][6] = 9'b110000000;
assign supra[6][7] = 9'b110100000;
assign supra[6][8] = 9'b110100000;
assign supra[6][9] = 9'b110100000;
assign supra[6][10] = 9'b110100000;
assign supra[6][11] = 9'b110100000;
assign supra[6][12] = 9'b110100000;
assign supra[6][13] = 9'b110000000;
assign supra[6][14] = 9'b110000000;
assign supra[6][15] = 9'b110100000;
assign supra[6][16] = 9'b110000000;
assign supra[6][17] = 9'b110100000;
assign supra[6][18] = 9'b110000000;
assign supra[7][1] = 9'b110000000;
assign supra[7][2] = 9'b110100000;
assign supra[7][3] = 9'b110000000;
assign supra[7][4] = 9'b110100000;
assign supra[7][5] = 9'b110000000;
assign supra[7][6] = 9'b110100000;
assign supra[7][7] = 9'b110100000;
assign supra[7][8] = 9'b110100000;
assign supra[7][9] = 9'b110100000;
assign supra[7][10] = 9'b110100000;
assign supra[7][11] = 9'b110100000;
assign supra[7][12] = 9'b110100000;
assign supra[7][13] = 9'b110100000;
assign supra[7][14] = 9'b110000000;
assign supra[7][15] = 9'b110100000;
assign supra[7][16] = 9'b110000000;
assign supra[7][17] = 9'b110100000;
assign supra[7][18] = 9'b110100000;
assign supra[8][1] = 9'b110100000;
assign supra[8][2] = 9'b110000000;
assign supra[8][3] = 9'b110100000;
assign supra[8][4] = 9'b110100000;
assign supra[8][5] = 9'b110000000;
assign supra[8][6] = 9'b110100000;
assign supra[8][7] = 9'b110100000;
assign supra[8][8] = 9'b110100000;
assign supra[8][9] = 9'b110100000;
assign supra[8][10] = 9'b110100000;
assign supra[8][11] = 9'b110100000;
assign supra[8][12] = 9'b110100000;
assign supra[8][13] = 9'b110100000;
assign supra[8][14] = 9'b110000000;
assign supra[8][15] = 9'b110100000;
assign supra[8][16] = 9'b110100000;
assign supra[8][17] = 9'b110000000;
assign supra[8][18] = 9'b110100000;
assign supra[9][1] = 9'b110100000;
assign supra[9][2] = 9'b110000000;
assign supra[9][3] = 9'b110100000;
assign supra[9][4] = 9'b110000000;
assign supra[9][5] = 9'b110000000;
assign supra[9][6] = 9'b110100000;
assign supra[9][7] = 9'b110100000;
assign supra[9][8] = 9'b110100000;
assign supra[9][9] = 9'b110100000;
assign supra[9][10] = 9'b110100000;
assign supra[9][11] = 9'b110100000;
assign supra[9][12] = 9'b110100000;
assign supra[9][13] = 9'b110100000;
assign supra[9][14] = 9'b110000000;
assign supra[9][15] = 9'b110000000;
assign supra[9][16] = 9'b110100000;
assign supra[9][17] = 9'b110000000;
assign supra[9][18] = 9'b110100000;
assign supra[10][1] = 9'b110100000;
assign supra[10][2] = 9'b110000000;
assign supra[10][3] = 9'b110100000;
assign supra[10][4] = 9'b110000000;
assign supra[10][5] = 9'b110000000;
assign supra[10][6] = 9'b110100000;
assign supra[10][7] = 9'b110100000;
assign supra[10][8] = 9'b110100000;
assign supra[10][9] = 9'b110100000;
assign supra[10][10] = 9'b110100000;
assign supra[10][11] = 9'b110100000;
assign supra[10][12] = 9'b110100000;
assign supra[10][13] = 9'b110100000;
assign supra[10][14] = 9'b110000000;
assign supra[10][15] = 9'b110000000;
assign supra[10][16] = 9'b110100000;
assign supra[10][17] = 9'b110000000;
assign supra[10][18] = 9'b110100000;
assign supra[11][1] = 9'b110100000;
assign supra[11][2] = 9'b110000000;
assign supra[11][3] = 9'b110100000;
assign supra[11][4] = 9'b110000000;
assign supra[11][5] = 9'b110000000;
assign supra[11][6] = 9'b110100000;
assign supra[11][7] = 9'b110100000;
assign supra[11][8] = 9'b110100000;
assign supra[11][9] = 9'b110100000;
assign supra[11][10] = 9'b110100000;
assign supra[11][11] = 9'b110100000;
assign supra[11][12] = 9'b110100000;
assign supra[11][13] = 9'b110100000;
assign supra[11][14] = 9'b110000000;
assign supra[11][15] = 9'b110000000;
assign supra[11][16] = 9'b110100000;
assign supra[11][17] = 9'b110000000;
assign supra[11][18] = 9'b110100000;
assign supra[12][1] = 9'b110100000;
assign supra[12][2] = 9'b110000000;
assign supra[12][3] = 9'b110100000;
assign supra[12][4] = 9'b110000000;
assign supra[12][5] = 9'b110000000;
assign supra[12][6] = 9'b110100000;
assign supra[12][7] = 9'b110100000;
assign supra[12][8] = 9'b110100000;
assign supra[12][9] = 9'b110100000;
assign supra[12][10] = 9'b110100000;
assign supra[12][11] = 9'b110100000;
assign supra[12][12] = 9'b110100000;
assign supra[12][13] = 9'b110100000;
assign supra[12][14] = 9'b110000000;
assign supra[12][15] = 9'b110000000;
assign supra[12][16] = 9'b110100000;
assign supra[12][17] = 9'b110000000;
assign supra[12][18] = 9'b110100000;
assign supra[13][1] = 9'b110100000;
assign supra[13][2] = 9'b110000000;
assign supra[13][3] = 9'b110100000;
assign supra[13][4] = 9'b110000000;
assign supra[13][5] = 9'b110000000;
assign supra[13][6] = 9'b110100000;
assign supra[13][7] = 9'b110100000;
assign supra[13][8] = 9'b110100000;
assign supra[13][9] = 9'b110100000;
assign supra[13][10] = 9'b110100000;
assign supra[13][11] = 9'b110100000;
assign supra[13][12] = 9'b110100000;
assign supra[13][13] = 9'b110100000;
assign supra[13][14] = 9'b110000000;
assign supra[13][15] = 9'b110000000;
assign supra[13][16] = 9'b110100000;
assign supra[13][17] = 9'b110000000;
assign supra[13][18] = 9'b110100000;
assign supra[13][19] = 9'b110000000;
assign supra[14][1] = 9'b110100000;
assign supra[14][2] = 9'b110000000;
assign supra[14][3] = 9'b110100000;
assign supra[14][4] = 9'b110000000;
assign supra[14][5] = 9'b110100000;
assign supra[14][6] = 9'b110100000;
assign supra[14][7] = 9'b110100000;
assign supra[14][8] = 9'b110100000;
assign supra[14][9] = 9'b110100000;
assign supra[14][10] = 9'b110100000;
assign supra[14][11] = 9'b110100000;
assign supra[14][12] = 9'b110100000;
assign supra[14][13] = 9'b110100000;
assign supra[14][14] = 9'b110100000;
assign supra[14][15] = 9'b110000000;
assign supra[14][16] = 9'b110100000;
assign supra[14][17] = 9'b110000000;
assign supra[14][18] = 9'b110100000;
assign supra[14][19] = 9'b110000000;
assign supra[15][1] = 9'b110100000;
assign supra[15][2] = 9'b110000000;
assign supra[15][3] = 9'b110100000;
assign supra[15][4] = 9'b110100000;
assign supra[15][5] = 9'b110000000;
assign supra[15][6] = 9'b101100000;
assign supra[15][7] = 9'b101000000;
assign supra[15][8] = 9'b101000000;
assign supra[15][9] = 9'b101000000;
assign supra[15][10] = 9'b101000000;
assign supra[15][11] = 9'b101000000;
assign supra[15][12] = 9'b101000000;
assign supra[15][13] = 9'b101100000;
assign supra[15][14] = 9'b110000000;
assign supra[15][15] = 9'b110100000;
assign supra[15][16] = 9'b110100000;
assign supra[15][17] = 9'b110000000;
assign supra[15][18] = 9'b110100000;
assign supra[15][19] = 9'b110000000;
assign supra[16][1] = 9'b110100000;
assign supra[16][2] = 9'b110100000;
assign supra[16][3] = 9'b110000000;
assign supra[16][4] = 9'b101000000;
assign supra[16][5] = 9'b100000000;
assign supra[16][6] = 9'b100000000;
assign supra[16][7] = 9'b100000000;
assign supra[16][8] = 9'b100000000;
assign supra[16][9] = 9'b100000000;
assign supra[16][10] = 9'b100000000;
assign supra[16][11] = 9'b100000000;
assign supra[16][12] = 9'b100000000;
assign supra[16][13] = 9'b100000000;
assign supra[16][14] = 9'b100000000;
assign supra[16][15] = 9'b101000000;
assign supra[16][16] = 9'b110000000;
assign supra[16][17] = 9'b110100000;
assign supra[16][18] = 9'b110100000;
assign supra[16][19] = 9'b110000000;
assign supra[17][1] = 9'b110100000;
assign supra[17][2] = 9'b110000000;
assign supra[17][3] = 9'b100100000;
assign supra[17][4] = 9'b100000000;
assign supra[17][5] = 9'b100000000;
assign supra[17][6] = 9'b100000100;
assign supra[17][7] = 9'b100001001;
assign supra[17][8] = 9'b100001001;
assign supra[17][9] = 9'b100001010;
assign supra[17][10] = 9'b100001010;
assign supra[17][11] = 9'b100001001;
assign supra[17][12] = 9'b100001001;
assign supra[17][13] = 9'b100000101;
assign supra[17][14] = 9'b100000100;
assign supra[17][15] = 9'b100000000;
assign supra[17][16] = 9'b100100000;
assign supra[17][17] = 9'b110000000;
assign supra[17][18] = 9'b110100000;
assign supra[18][1] = 9'b111100000;
assign supra[18][2] = 9'b101000000;
assign supra[18][3] = 9'b100000100;
assign supra[18][4] = 9'b100001001;
assign supra[18][5] = 9'b100001010;
assign supra[18][6] = 9'b100001111;
assign supra[18][7] = 9'b100001111;
assign supra[18][8] = 9'b100001111;
assign supra[18][9] = 9'b100001111;
assign supra[18][10] = 9'b100001111;
assign supra[18][11] = 9'b100001111;
assign supra[18][12] = 9'b100001111;
assign supra[18][13] = 9'b100001111;
assign supra[18][14] = 9'b100001111;
assign supra[18][15] = 9'b100001111;
assign supra[18][16] = 9'b100000101;
assign supra[18][17] = 9'b101000000;
assign supra[18][18] = 9'b111100000;
assign supra[19][1] = 9'b111100000;
assign supra[19][2] = 9'b101100000;
assign supra[19][3] = 9'b100001111;
assign supra[19][4] = 9'b100001111;
assign supra[19][5] = 9'b100001111;
assign supra[19][6] = 9'b100001111;
assign supra[19][7] = 9'b100001111;
assign supra[19][8] = 9'b100001111;
assign supra[19][9] = 9'b100001111;
assign supra[19][10] = 9'b100001111;
assign supra[19][11] = 9'b100001111;
assign supra[19][12] = 9'b100001111;
assign supra[19][13] = 9'b100001111;
assign supra[19][14] = 9'b100001111;
assign supra[19][15] = 9'b100001111;
assign supra[19][16] = 9'b100001111;
assign supra[19][17] = 9'b101000000;
assign supra[19][18] = 9'b111100000;
assign supra[20][1] = 9'b110100000;
assign supra[20][2] = 9'b101100000;
assign supra[20][3] = 9'b100001011;
assign supra[20][4] = 9'b100001111;
assign supra[20][5] = 9'b100001111;
assign supra[20][6] = 9'b100001111;
assign supra[20][7] = 9'b100001111;
assign supra[20][8] = 9'b100001111;
assign supra[20][9] = 9'b100001111;
assign supra[20][10] = 9'b100001111;
assign supra[20][11] = 9'b100001011;
assign supra[20][12] = 9'b100001111;
assign supra[20][13] = 9'b100001111;
assign supra[20][14] = 9'b100001111;
assign supra[20][15] = 9'b100001111;
assign supra[20][16] = 9'b100001010;
assign supra[20][17] = 9'b101100000;
assign supra[20][18] = 9'b110100000;
assign supra[21][0] = 9'b110000000;
assign supra[21][1] = 9'b110000000;
assign supra[21][2] = 9'b101000101;
assign supra[21][3] = 9'b100100101;
assign supra[21][4] = 9'b100000110;
assign supra[21][5] = 9'b100001111;
assign supra[21][6] = 9'b100001111;
assign supra[21][7] = 9'b100001011;
assign supra[21][8] = 9'b100001010;
assign supra[21][9] = 9'b100001111;
assign supra[21][10] = 9'b100001111;
assign supra[21][11] = 9'b100001010;
assign supra[21][12] = 9'b100000101;
assign supra[21][13] = 9'b100000101;
assign supra[21][14] = 9'b100000101;
assign supra[21][15] = 9'b100000110;
assign supra[21][16] = 9'b100100101;
assign supra[21][17] = 9'b101000101;
assign supra[21][18] = 9'b110000000;
assign supra[21][19] = 9'b110000000;
assign supra[22][0] = 9'b110000000;
assign supra[22][1] = 9'b110100000;
assign supra[22][2] = 9'b100101001;
assign supra[22][3] = 9'b100100000;
assign supra[22][4] = 9'b100000001;
assign supra[22][5] = 9'b100001010;
assign supra[22][6] = 9'b100001010;
assign supra[22][7] = 9'b100000001;
assign supra[22][8] = 9'b100000001;
assign supra[22][9] = 9'b100001111;
assign supra[22][10] = 9'b100001111;
assign supra[22][11] = 9'b100000101;
assign supra[22][12] = 9'b100000001;
assign supra[22][13] = 9'b100000001;
assign supra[22][14] = 9'b100000001;
assign supra[22][15] = 9'b100000001;
assign supra[22][16] = 9'b100100000;
assign supra[22][17] = 9'b100101001;
assign supra[22][18] = 9'b110100000;
assign supra[22][19] = 9'b110000000;
assign supra[23][1] = 9'b110100000;
assign supra[23][2] = 9'b100101010;
assign supra[23][3] = 9'b101000101;
assign supra[23][4] = 9'b100001010;
assign supra[23][5] = 9'b100001111;
assign supra[23][6] = 9'b100001111;
assign supra[23][7] = 9'b100001111;
assign supra[23][8] = 9'b100001011;
assign supra[23][9] = 9'b100001111;
assign supra[23][10] = 9'b100001111;
assign supra[23][11] = 9'b100001011;
assign supra[23][12] = 9'b100001111;
assign supra[23][13] = 9'b100010011;
assign supra[23][14] = 9'b100010011;
assign supra[23][15] = 9'b100001111;
assign supra[23][16] = 9'b101000101;
assign supra[23][17] = 9'b100001010;
assign supra[23][18] = 9'b110100000;
assign supra[24][1] = 9'b110100000;
assign supra[24][2] = 9'b100001010;
assign supra[24][3] = 9'b100101001;
assign supra[24][4] = 9'b101100000;
assign supra[24][5] = 9'b100101001;
assign supra[24][6] = 9'b100100101;
assign supra[24][7] = 9'b101000101;
assign supra[24][8] = 9'b101000100;
assign supra[24][9] = 9'b101000100;
assign supra[24][10] = 9'b101000100;
assign supra[24][11] = 9'b101000100;
assign supra[24][12] = 9'b101000101;
assign supra[24][13] = 9'b100100101;
assign supra[24][14] = 9'b100101001;
assign supra[24][15] = 9'b101100000;
assign supra[24][16] = 9'b100101001;
assign supra[24][17] = 9'b100001010;
assign supra[24][18] = 9'b110100000;
assign supra[25][1] = 9'b110100000;
assign supra[25][2] = 9'b100101001;
assign supra[25][3] = 9'b100001111;
assign supra[25][4] = 9'b110000000;
assign supra[25][5] = 9'b110100000;
assign supra[25][6] = 9'b110100000;
assign supra[25][7] = 9'b110100000;
assign supra[25][8] = 9'b110100000;
assign supra[25][9] = 9'b110100000;
assign supra[25][10] = 9'b110100000;
assign supra[25][11] = 9'b110100000;
assign supra[25][12] = 9'b110100000;
assign supra[25][13] = 9'b110100000;
assign supra[25][14] = 9'b110100000;
assign supra[25][15] = 9'b110000000;
assign supra[25][16] = 9'b100001111;
assign supra[25][17] = 9'b100101010;
assign supra[25][18] = 9'b110100000;
assign supra[26][1] = 9'b110100000;
assign supra[26][2] = 9'b100101001;
assign supra[26][3] = 9'b100001111;
assign supra[26][4] = 9'b101100000;
assign supra[26][5] = 9'b110100000;
assign supra[26][6] = 9'b110100000;
assign supra[26][7] = 9'b110100000;
assign supra[26][8] = 9'b110100000;
assign supra[26][9] = 9'b110100000;
assign supra[26][10] = 9'b110100000;
assign supra[26][11] = 9'b110100000;
assign supra[26][12] = 9'b110100000;
assign supra[26][13] = 9'b110100000;
assign supra[26][14] = 9'b110100000;
assign supra[26][15] = 9'b101100000;
assign supra[26][16] = 9'b100001111;
assign supra[26][17] = 9'b100101001;
assign supra[26][18] = 9'b110100000;
assign supra[27][1] = 9'b110100000;
assign supra[27][2] = 9'b100101001;
assign supra[27][3] = 9'b100001111;
assign supra[27][4] = 9'b101100000;
assign supra[27][5] = 9'b110100000;
assign supra[27][6] = 9'b110100000;
assign supra[27][7] = 9'b110100000;
assign supra[27][8] = 9'b110100000;
assign supra[27][9] = 9'b110100000;
assign supra[27][10] = 9'b110100000;
assign supra[27][11] = 9'b110100000;
assign supra[27][12] = 9'b110100000;
assign supra[27][13] = 9'b110100000;
assign supra[27][14] = 9'b110100000;
assign supra[27][15] = 9'b101100000;
assign supra[27][16] = 9'b100001111;
assign supra[27][17] = 9'b100101001;
assign supra[27][18] = 9'b110100000;
assign supra[28][1] = 9'b110100000;
assign supra[28][2] = 9'b100101001;
assign supra[28][3] = 9'b100001111;
assign supra[28][4] = 9'b101100100;
assign supra[28][5] = 9'b110100000;
assign supra[28][6] = 9'b110100000;
assign supra[28][7] = 9'b110100000;
assign supra[28][8] = 9'b110100000;
assign supra[28][9] = 9'b110100000;
assign supra[28][10] = 9'b110100000;
assign supra[28][11] = 9'b110100000;
assign supra[28][12] = 9'b110100000;
assign supra[28][13] = 9'b110100000;
assign supra[28][14] = 9'b110100000;
assign supra[28][15] = 9'b101100000;
assign supra[28][16] = 9'b100001111;
assign supra[28][17] = 9'b100101001;
assign supra[28][18] = 9'b110100000;
assign supra[29][1] = 9'b110100000;
assign supra[29][2] = 9'b100100101;
assign supra[29][3] = 9'b100001111;
assign supra[29][4] = 9'b101100000;
assign supra[29][5] = 9'b110100000;
assign supra[29][6] = 9'b110100000;
assign supra[29][7] = 9'b110100000;
assign supra[29][8] = 9'b110100000;
assign supra[29][9] = 9'b110100000;
assign supra[29][10] = 9'b110100000;
assign supra[29][11] = 9'b110100000;
assign supra[29][12] = 9'b110100000;
assign supra[29][13] = 9'b110100000;
assign supra[29][14] = 9'b110100000;
assign supra[29][15] = 9'b101100000;
assign supra[29][16] = 9'b100001111;
assign supra[29][17] = 9'b100101001;
assign supra[29][18] = 9'b110100000;
assign supra[30][1] = 9'b110100000;
assign supra[30][2] = 9'b100100101;
assign supra[30][3] = 9'b100001011;
assign supra[30][4] = 9'b101100000;
assign supra[30][5] = 9'b110100000;
assign supra[30][6] = 9'b110100000;
assign supra[30][7] = 9'b110100000;
assign supra[30][8] = 9'b110100000;
assign supra[30][9] = 9'b110100000;
assign supra[30][10] = 9'b110100000;
assign supra[30][11] = 9'b110100000;
assign supra[30][12] = 9'b110100000;
assign supra[30][13] = 9'b110100000;
assign supra[30][14] = 9'b110100000;
assign supra[30][15] = 9'b101100000;
assign supra[30][16] = 9'b100001011;
assign supra[30][17] = 9'b100100101;
assign supra[30][18] = 9'b110100000;
assign supra[31][1] = 9'b110100000;
assign supra[31][2] = 9'b100100101;
assign supra[31][3] = 9'b100000101;
assign supra[31][4] = 9'b110000000;
assign supra[31][5] = 9'b110000000;
assign supra[31][6] = 9'b110100000;
assign supra[31][7] = 9'b110100000;
assign supra[31][8] = 9'b110100000;
assign supra[31][9] = 9'b110100000;
assign supra[31][10] = 9'b110100000;
assign supra[31][11] = 9'b110100000;
assign supra[31][12] = 9'b110100000;
assign supra[31][13] = 9'b110100000;
assign supra[31][14] = 9'b110000000;
assign supra[31][15] = 9'b110000000;
assign supra[31][16] = 9'b100000101;
assign supra[31][17] = 9'b100100101;
assign supra[31][18] = 9'b110100000;
assign supra[32][1] = 9'b110100000;
assign supra[32][2] = 9'b100100101;
assign supra[32][3] = 9'b100000001;
assign supra[32][4] = 9'b110000000;
assign supra[32][5] = 9'b110000000;
assign supra[32][6] = 9'b110100000;
assign supra[32][7] = 9'b110100000;
assign supra[32][8] = 9'b110100000;
assign supra[32][9] = 9'b110100000;
assign supra[32][10] = 9'b110100000;
assign supra[32][11] = 9'b110100000;
assign supra[32][12] = 9'b110100000;
assign supra[32][13] = 9'b110100000;
assign supra[32][14] = 9'b110000000;
assign supra[32][15] = 9'b110000000;
assign supra[32][16] = 9'b100000001;
assign supra[32][17] = 9'b100100101;
assign supra[32][18] = 9'b110100000;
assign supra[33][1] = 9'b110100000;
assign supra[33][2] = 9'b100100101;
assign supra[33][3] = 9'b100000001;
assign supra[33][4] = 9'b110100000;
assign supra[33][5] = 9'b110000000;
assign supra[33][6] = 9'b110100000;
assign supra[33][7] = 9'b110100000;
assign supra[33][8] = 9'b110100000;
assign supra[33][9] = 9'b110100000;
assign supra[33][10] = 9'b110100000;
assign supra[33][11] = 9'b110100000;
assign supra[33][12] = 9'b110100000;
assign supra[33][13] = 9'b110100000;
assign supra[33][14] = 9'b110000000;
assign supra[33][15] = 9'b110100000;
assign supra[33][16] = 9'b100100001;
assign supra[33][17] = 9'b100101001;
assign supra[33][18] = 9'b110100000;
assign supra[34][0] = 9'b101100100;
assign supra[34][1] = 9'b110100000;
assign supra[34][2] = 9'b100100101;
assign supra[34][3] = 9'b101000101;
assign supra[34][4] = 9'b111100000;
assign supra[34][5] = 9'b110000000;
assign supra[34][6] = 9'b110000000;
assign supra[34][7] = 9'b110000000;
assign supra[34][8] = 9'b110000000;
assign supra[34][9] = 9'b110000000;
assign supra[34][10] = 9'b110000000;
assign supra[34][11] = 9'b110000000;
assign supra[34][12] = 9'b110000000;
assign supra[34][13] = 9'b110000000;
assign supra[34][14] = 9'b110000000;
assign supra[34][15] = 9'b110100000;
assign supra[34][16] = 9'b101000101;
assign supra[34][17] = 9'b100100101;
assign supra[34][18] = 9'b110100000;
assign supra[34][19] = 9'b101100100;
assign supra[35][0] = 9'b101100100;
assign supra[35][1] = 9'b110100000;
assign supra[35][2] = 9'b110000000;
assign supra[35][3] = 9'b110000000;
assign supra[35][4] = 9'b110000000;
assign supra[35][5] = 9'b100001001;
assign supra[35][6] = 9'b100001010;
assign supra[35][7] = 9'b100001010;
assign supra[35][8] = 9'b100001010;
assign supra[35][9] = 9'b100101101;
assign supra[35][10] = 9'b100101101;
assign supra[35][11] = 9'b100001010;
assign supra[35][12] = 9'b100001010;
assign supra[35][13] = 9'b100001010;
assign supra[35][14] = 9'b100001001;
assign supra[35][15] = 9'b101100000;
assign supra[35][16] = 9'b110000000;
assign supra[35][17] = 9'b110000000;
assign supra[35][18] = 9'b110100000;
assign supra[35][19] = 9'b101100100;
assign supra[36][0] = 9'b110000000;
assign supra[36][1] = 9'b110000000;
assign supra[36][2] = 9'b110100000;
assign supra[36][3] = 9'b110100000;
assign supra[36][4] = 9'b100100100;
assign supra[36][5] = 9'b100001111;
assign supra[36][6] = 9'b100001111;
assign supra[36][7] = 9'b100001111;
assign supra[36][8] = 9'b100001111;
assign supra[36][9] = 9'b100001111;
assign supra[36][10] = 9'b100001111;
assign supra[36][11] = 9'b100001111;
assign supra[36][12] = 9'b100001111;
assign supra[36][13] = 9'b100001111;
assign supra[36][14] = 9'b100001111;
assign supra[36][15] = 9'b100100101;
assign supra[36][16] = 9'b110100000;
assign supra[36][17] = 9'b110100000;
assign supra[36][18] = 9'b110000000;
assign supra[36][19] = 9'b110000000;
assign supra[37][0] = 9'b110000000;
assign supra[37][1] = 9'b110000000;
assign supra[37][2] = 9'b110100000;
assign supra[37][3] = 9'b110100000;
assign supra[37][4] = 9'b100100101;
assign supra[37][5] = 9'b100001111;
assign supra[37][6] = 9'b100001111;
assign supra[37][7] = 9'b100001111;
assign supra[37][8] = 9'b100001111;
assign supra[37][9] = 9'b100001111;
assign supra[37][10] = 9'b100001111;
assign supra[37][11] = 9'b100001111;
assign supra[37][12] = 9'b100001111;
assign supra[37][13] = 9'b100001111;
assign supra[37][14] = 9'b100001111;
assign supra[37][15] = 9'b100101001;
assign supra[37][16] = 9'b110100000;
assign supra[37][17] = 9'b110100000;
assign supra[37][18] = 9'b110000000;
assign supra[37][19] = 9'b110000000;
assign supra[38][0] = 9'b110000000;
assign supra[38][1] = 9'b110000000;
assign supra[38][2] = 9'b110100000;
assign supra[38][3] = 9'b110000000;
assign supra[38][4] = 9'b100001010;
assign supra[38][5] = 9'b100001111;
assign supra[38][6] = 9'b100001111;
assign supra[38][7] = 9'b100001111;
assign supra[38][8] = 9'b100001111;
assign supra[38][9] = 9'b100001111;
assign supra[38][10] = 9'b100001111;
assign supra[38][11] = 9'b100001111;
assign supra[38][12] = 9'b100001111;
assign supra[38][13] = 9'b100001111;
assign supra[38][14] = 9'b100001111;
assign supra[38][15] = 9'b100001010;
assign supra[38][16] = 9'b110000000;
assign supra[38][17] = 9'b110100000;
assign supra[38][18] = 9'b110000000;
assign supra[38][19] = 9'b110000000;
assign supra[39][0] = 9'b110000000;
assign supra[39][1] = 9'b110000000;
assign supra[39][2] = 9'b110100000;
assign supra[39][3] = 9'b110000000;
assign supra[39][4] = 9'b100001011;
assign supra[39][5] = 9'b100001111;
assign supra[39][6] = 9'b100001111;
assign supra[39][7] = 9'b100001111;
assign supra[39][8] = 9'b100001111;
assign supra[39][9] = 9'b100001111;
assign supra[39][10] = 9'b100001111;
assign supra[39][11] = 9'b100001111;
assign supra[39][12] = 9'b100001111;
assign supra[39][13] = 9'b100001111;
assign supra[39][14] = 9'b100001111;
assign supra[39][15] = 9'b100001011;
assign supra[39][16] = 9'b110000000;
assign supra[39][17] = 9'b110100000;
assign supra[39][18] = 9'b110000000;
assign supra[39][19] = 9'b110000000;
assign supra[40][0] = 9'b110000000;
assign supra[40][1] = 9'b110000000;
assign supra[40][2] = 9'b110100000;
assign supra[40][3] = 9'b101100000;
assign supra[40][4] = 9'b100001111;
assign supra[40][5] = 9'b100001111;
assign supra[40][6] = 9'b100001111;
assign supra[40][7] = 9'b100001111;
assign supra[40][8] = 9'b100001111;
assign supra[40][9] = 9'b100001111;
assign supra[40][10] = 9'b100001111;
assign supra[40][11] = 9'b100001111;
assign supra[40][12] = 9'b100001111;
assign supra[40][13] = 9'b100001111;
assign supra[40][14] = 9'b100001111;
assign supra[40][15] = 9'b100001111;
assign supra[40][16] = 9'b101100000;
assign supra[40][17] = 9'b110100000;
assign supra[40][18] = 9'b110000000;
assign supra[40][19] = 9'b110000000;
assign supra[41][0] = 9'b110100000;
assign supra[41][1] = 9'b110000000;
assign supra[41][2] = 9'b110000000;
assign supra[41][3] = 9'b101100000;
assign supra[41][4] = 9'b100001111;
assign supra[41][5] = 9'b100001111;
assign supra[41][6] = 9'b100001111;
assign supra[41][7] = 9'b100001111;
assign supra[41][8] = 9'b100001111;
assign supra[41][9] = 9'b100001111;
assign supra[41][10] = 9'b100001111;
assign supra[41][11] = 9'b100001111;
assign supra[41][12] = 9'b100001111;
assign supra[41][13] = 9'b100001111;
assign supra[41][14] = 9'b100001111;
assign supra[41][15] = 9'b100001111;
assign supra[41][16] = 9'b101100000;
assign supra[41][17] = 9'b110100000;
assign supra[41][18] = 9'b110000000;
assign supra[41][19] = 9'b110100000;
assign supra[42][0] = 9'b110100000;
assign supra[42][1] = 9'b110000000;
assign supra[42][2] = 9'b110000000;
assign supra[42][3] = 9'b110000000;
assign supra[42][4] = 9'b100001001;
assign supra[42][5] = 9'b100001111;
assign supra[42][6] = 9'b100001111;
assign supra[42][7] = 9'b100001111;
assign supra[42][8] = 9'b100001111;
assign supra[42][9] = 9'b100001111;
assign supra[42][10] = 9'b100001111;
assign supra[42][11] = 9'b100001111;
assign supra[42][12] = 9'b100001111;
assign supra[42][13] = 9'b100001111;
assign supra[42][14] = 9'b100001111;
assign supra[42][15] = 9'b100001001;
assign supra[42][16] = 9'b110000000;
assign supra[42][17] = 9'b110000000;
assign supra[42][18] = 9'b110000000;
assign supra[42][19] = 9'b110100000;
assign supra[43][1] = 9'b110000000;
assign supra[43][2] = 9'b110000000;
assign supra[43][3] = 9'b110100000;
assign supra[43][4] = 9'b101100000;
assign supra[43][5] = 9'b100001001;
assign supra[43][6] = 9'b100001111;
assign supra[43][7] = 9'b100001111;
assign supra[43][8] = 9'b100001111;
assign supra[43][9] = 9'b100001111;
assign supra[43][10] = 9'b100001111;
assign supra[43][11] = 9'b100001111;
assign supra[43][12] = 9'b100001111;
assign supra[43][13] = 9'b100001111;
assign supra[43][14] = 9'b100001001;
assign supra[43][15] = 9'b101100000;
assign supra[43][16] = 9'b110100000;
assign supra[43][17] = 9'b110000000;
assign supra[43][18] = 9'b110000000;
assign supra[44][1] = 9'b110000000;
assign supra[44][2] = 9'b110000000;
assign supra[44][3] = 9'b110000000;
assign supra[44][4] = 9'b110100000;
assign supra[44][5] = 9'b110000000;
assign supra[44][6] = 9'b101100000;
assign supra[44][7] = 9'b101000000;
assign supra[44][8] = 9'b100100101;
assign supra[44][9] = 9'b100100101;
assign supra[44][10] = 9'b100100101;
assign supra[44][11] = 9'b100100101;
assign supra[44][12] = 9'b101000100;
assign supra[44][13] = 9'b101100000;
assign supra[44][14] = 9'b110000000;
assign supra[44][15] = 9'b110100000;
assign supra[44][16] = 9'b110000000;
assign supra[44][17] = 9'b110000000;
assign supra[44][18] = 9'b110000000;
assign supra[45][1] = 9'b110000000;
assign supra[45][2] = 9'b110000000;
assign supra[45][3] = 9'b110000000;
assign supra[45][4] = 9'b110000000;
assign supra[45][5] = 9'b110100000;
assign supra[45][6] = 9'b110100000;
assign supra[45][7] = 9'b110100000;
assign supra[45][8] = 9'b110100000;
assign supra[45][9] = 9'b110100000;
assign supra[45][10] = 9'b110100000;
assign supra[45][11] = 9'b110100000;
assign supra[45][12] = 9'b110100000;
assign supra[45][13] = 9'b110100000;
assign supra[45][14] = 9'b110100000;
assign supra[45][15] = 9'b110000000;
assign supra[45][16] = 9'b110000000;
assign supra[45][17] = 9'b110000000;
assign supra[45][18] = 9'b110000000;
assign supra[46][2] = 9'b110000100;
assign supra[46][3] = 9'b110101101;
assign supra[46][4] = 9'b110101101;
assign supra[46][5] = 9'b110101101;
assign supra[46][6] = 9'b110101101;
assign supra[46][7] = 9'b110101101;
assign supra[46][8] = 9'b110101101;
assign supra[46][9] = 9'b110101101;
assign supra[46][10] = 9'b110101101;
assign supra[46][11] = 9'b110101101;
assign supra[46][12] = 9'b110101101;
assign supra[46][13] = 9'b110101101;
assign supra[46][14] = 9'b110101101;
assign supra[46][15] = 9'b110101101;
assign supra[46][16] = 9'b110101101;
assign supra[46][17] = 9'b110000100;
assign supra[47][2] = 9'b110000100;
assign supra[47][3] = 9'b111111111;
assign supra[47][4] = 9'b111111111;
assign supra[47][5] = 9'b111111111;
assign supra[47][6] = 9'b111111111;
assign supra[47][7] = 9'b111111111;
assign supra[47][8] = 9'b111111111;
assign supra[47][9] = 9'b111111111;
assign supra[47][10] = 9'b111111111;
assign supra[47][11] = 9'b111111111;
assign supra[47][12] = 9'b111111111;
assign supra[47][13] = 9'b111111111;
assign supra[47][14] = 9'b111111111;
assign supra[47][15] = 9'b111111111;
assign supra[47][16] = 9'b111111111;
assign supra[47][17] = 9'b110000100;
assign supra[48][2] = 9'b110001101;
assign supra[48][3] = 9'b111110110;
assign supra[48][4] = 9'b111110110;
assign supra[48][5] = 9'b111110010;
assign supra[48][6] = 9'b111110110;
assign supra[48][7] = 9'b111110110;
assign supra[48][8] = 9'b111110110;
assign supra[48][9] = 9'b111110110;
assign supra[48][10] = 9'b111110110;
assign supra[48][11] = 9'b111110110;
assign supra[48][12] = 9'b111110110;
assign supra[48][13] = 9'b111110110;
assign supra[48][14] = 9'b111110010;
assign supra[48][15] = 9'b111110110;
assign supra[48][16] = 9'b111110110;
assign supra[48][17] = 9'b110001101;
assign supra[49][4] = 9'b110000000;
assign supra[49][5] = 9'b110000000;
assign supra[49][6] = 9'b110000000;
assign supra[49][7] = 9'b110000000;
assign supra[49][8] = 9'b110000000;
assign supra[49][9] = 9'b110000000;
assign supra[49][10] = 9'b110000000;
assign supra[49][11] = 9'b110000000;
assign supra[49][12] = 9'b110000000;
assign supra[49][13] = 9'b110000000;
assign supra[49][14] = 9'b110000000;
assign supra[49][15] = 9'b110000000;
//Total de Lineas = 900
endmodule

