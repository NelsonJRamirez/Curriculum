`timescale 1ns / 1ps
module reset_logo (
input enable,
input clock,
input [9:0] posx, posy,
input [9:0] hcount,
input [9:0] vcount,
output reg[2:0] red,
output reg[2:0] green,
output reg[1:0] blue,
output reg data);

always @(posedge clock)
begin
	if(enable)
	begin
		if(hcount >= posx & hcount < posx + RESOLUCION_X & vcount >= posy & vcount < posy + RESOLUCION_Y)
		begin
			if (reset_logo[vcount - posy][hcount - posx][8] == 1'b1)
			begin
				red   <= reset_logo[vcount- posy][hcount- posx][7:5];
				green <= reset_logo[vcount- posy][hcount- posx][4:2];
            blue 	<= reset_logo[vcount- posy][hcount- posx][1:0];
				data  <= 1'b1;
			end
			else
				data <= 0;
			end
		else
		data <= 0;
	end
end

parameter RESOLUCION_X = 40;
parameter RESOLUCION_Y = 40;
wire [8:0] reset_logo[RESOLUCION_Y - 1'b1 : 0][RESOLUCION_X - 1'b1 : 0];
assign reset_logo[0][15] = 9'b100100100;
assign reset_logo[0][16] = 9'b100100100;
assign reset_logo[0][17] = 9'b101001000;
assign reset_logo[0][18] = 9'b101001000;
assign reset_logo[0][19] = 9'b101001001;
assign reset_logo[0][20] = 9'b101001001;
assign reset_logo[0][21] = 9'b101001001;
assign reset_logo[0][22] = 9'b101001001;
assign reset_logo[0][23] = 9'b101001001;
assign reset_logo[0][24] = 9'b101001001;
assign reset_logo[1][12] = 9'b100100100;
assign reset_logo[1][13] = 9'b101001000;
assign reset_logo[1][14] = 9'b101001000;
assign reset_logo[1][15] = 9'b101001001;
assign reset_logo[1][16] = 9'b101001001;
assign reset_logo[1][17] = 9'b101001001;
assign reset_logo[1][18] = 9'b101001001;
assign reset_logo[1][19] = 9'b101101101;
assign reset_logo[1][20] = 9'b101101101;
assign reset_logo[1][21] = 9'b101001001;
assign reset_logo[1][22] = 9'b101001001;
assign reset_logo[1][23] = 9'b101101101;
assign reset_logo[1][24] = 9'b101101101;
assign reset_logo[1][25] = 9'b101101101;
assign reset_logo[1][26] = 9'b101101101;
assign reset_logo[1][27] = 9'b101001001;
assign reset_logo[2][10] = 9'b100100100;
assign reset_logo[2][11] = 9'b100100100;
assign reset_logo[2][12] = 9'b101001000;
assign reset_logo[2][13] = 9'b101001000;
assign reset_logo[2][14] = 9'b101001001;
assign reset_logo[2][15] = 9'b101001001;
assign reset_logo[2][16] = 9'b101101101;
assign reset_logo[2][17] = 9'b101101101;
assign reset_logo[2][18] = 9'b101101101;
assign reset_logo[2][19] = 9'b101101101;
assign reset_logo[2][20] = 9'b101101101;
assign reset_logo[2][21] = 9'b101101101;
assign reset_logo[2][22] = 9'b101101101;
assign reset_logo[2][23] = 9'b101101101;
assign reset_logo[2][24] = 9'b101101101;
assign reset_logo[2][25] = 9'b101101101;
assign reset_logo[2][26] = 9'b101101101;
assign reset_logo[2][27] = 9'b101101101;
assign reset_logo[2][28] = 9'b101101101;
assign reset_logo[2][29] = 9'b101001001;
assign reset_logo[3][8] = 9'b100100100;
assign reset_logo[3][9] = 9'b100100100;
assign reset_logo[3][10] = 9'b100100100;
assign reset_logo[3][11] = 9'b101001000;
assign reset_logo[3][12] = 9'b101001001;
assign reset_logo[3][13] = 9'b101001001;
assign reset_logo[3][14] = 9'b101101101;
assign reset_logo[3][15] = 9'b101101101;
assign reset_logo[3][16] = 9'b101101101;
assign reset_logo[3][17] = 9'b101101101;
assign reset_logo[3][18] = 9'b101101101;
assign reset_logo[3][19] = 9'b110010001;
assign reset_logo[3][20] = 9'b110001101;
assign reset_logo[3][21] = 9'b101101101;
assign reset_logo[3][22] = 9'b101101101;
assign reset_logo[3][23] = 9'b101001001;
assign reset_logo[3][24] = 9'b101101101;
assign reset_logo[3][25] = 9'b101101101;
assign reset_logo[3][26] = 9'b101101101;
assign reset_logo[3][27] = 9'b101101101;
assign reset_logo[3][28] = 9'b101101101;
assign reset_logo[3][29] = 9'b101101101;
assign reset_logo[3][30] = 9'b101101101;
assign reset_logo[3][31] = 9'b101001001;
assign reset_logo[4][7] = 9'b100100100;
assign reset_logo[4][8] = 9'b100100100;
assign reset_logo[4][9] = 9'b100100100;
assign reset_logo[4][10] = 9'b101001001;
assign reset_logo[4][11] = 9'b101001001;
assign reset_logo[4][12] = 9'b101001001;
assign reset_logo[4][13] = 9'b101101101;
assign reset_logo[4][14] = 9'b101101101;
assign reset_logo[4][15] = 9'b101101101;
assign reset_logo[4][16] = 9'b101101101;
assign reset_logo[4][17] = 9'b110010001;
assign reset_logo[4][18] = 9'b110010001;
assign reset_logo[4][19] = 9'b110010001;
assign reset_logo[4][20] = 9'b110010001;
assign reset_logo[4][21] = 9'b101110001;
assign reset_logo[4][22] = 9'b101101101;
assign reset_logo[4][23] = 9'b101101101;
assign reset_logo[4][24] = 9'b101001001;
assign reset_logo[4][25] = 9'b101101001;
assign reset_logo[4][26] = 9'b101101101;
assign reset_logo[4][27] = 9'b101101101;
assign reset_logo[4][28] = 9'b101101101;
assign reset_logo[4][29] = 9'b101101101;
assign reset_logo[4][30] = 9'b101101101;
assign reset_logo[4][31] = 9'b101101101;
assign reset_logo[4][32] = 9'b101001001;
assign reset_logo[5][6] = 9'b100100100;
assign reset_logo[5][7] = 9'b100100100;
assign reset_logo[5][8] = 9'b100100100;
assign reset_logo[5][9] = 9'b101001001;
assign reset_logo[5][10] = 9'b101001001;
assign reset_logo[5][11] = 9'b101001001;
assign reset_logo[5][12] = 9'b101101101;
assign reset_logo[5][13] = 9'b101101101;
assign reset_logo[5][14] = 9'b101101101;
assign reset_logo[5][15] = 9'b110010001;
assign reset_logo[5][16] = 9'b110001101;
assign reset_logo[5][17] = 9'b110101101;
assign reset_logo[5][18] = 9'b111101001;
assign reset_logo[5][19] = 9'b111101001;
assign reset_logo[5][20] = 9'b111101001;
assign reset_logo[5][21] = 9'b111101001;
assign reset_logo[5][22] = 9'b110101101;
assign reset_logo[5][23] = 9'b110001101;
assign reset_logo[5][24] = 9'b101101101;
assign reset_logo[5][25] = 9'b101101101;
assign reset_logo[5][26] = 9'b101001101;
assign reset_logo[5][27] = 9'b101101001;
assign reset_logo[5][28] = 9'b101101101;
assign reset_logo[5][29] = 9'b101101101;
assign reset_logo[5][30] = 9'b101101101;
assign reset_logo[5][31] = 9'b101001001;
assign reset_logo[5][32] = 9'b101101101;
assign reset_logo[5][33] = 9'b101001001;
assign reset_logo[6][5] = 9'b100100100;
assign reset_logo[6][6] = 9'b100100100;
assign reset_logo[6][7] = 9'b101001000;
assign reset_logo[6][8] = 9'b101001001;
assign reset_logo[6][9] = 9'b101001001;
assign reset_logo[6][10] = 9'b101101001;
assign reset_logo[6][11] = 9'b101101101;
assign reset_logo[6][12] = 9'b101101101;
assign reset_logo[6][13] = 9'b110001101;
assign reset_logo[6][14] = 9'b111101101;
assign reset_logo[6][15] = 9'b111101000;
assign reset_logo[6][16] = 9'b111101000;
assign reset_logo[6][17] = 9'b111101000;
assign reset_logo[6][18] = 9'b111101000;
assign reset_logo[6][19] = 9'b111101000;
assign reset_logo[6][20] = 9'b111101000;
assign reset_logo[6][21] = 9'b111101000;
assign reset_logo[6][22] = 9'b111101000;
assign reset_logo[6][23] = 9'b111101000;
assign reset_logo[6][24] = 9'b111101001;
assign reset_logo[6][25] = 9'b111101001;
assign reset_logo[6][26] = 9'b110001101;
assign reset_logo[6][27] = 9'b101101101;
assign reset_logo[6][28] = 9'b101001001;
assign reset_logo[6][29] = 9'b101101001;
assign reset_logo[6][30] = 9'b101101101;
assign reset_logo[6][31] = 9'b101101101;
assign reset_logo[6][32] = 9'b101001001;
assign reset_logo[6][33] = 9'b101101101;
assign reset_logo[6][34] = 9'b101001001;
assign reset_logo[7][4] = 9'b100100100;
assign reset_logo[7][5] = 9'b100100100;
assign reset_logo[7][6] = 9'b101001000;
assign reset_logo[7][7] = 9'b101001001;
assign reset_logo[7][8] = 9'b101001001;
assign reset_logo[7][9] = 9'b101101001;
assign reset_logo[7][10] = 9'b101101101;
assign reset_logo[7][11] = 9'b110010001;
assign reset_logo[7][12] = 9'b111101101;
assign reset_logo[7][13] = 9'b111101000;
assign reset_logo[7][14] = 9'b111100100;
assign reset_logo[7][15] = 9'b111100100;
assign reset_logo[7][16] = 9'b111101000;
assign reset_logo[7][17] = 9'b111101000;
assign reset_logo[7][18] = 9'b111101001;
assign reset_logo[7][19] = 9'b111101101;
assign reset_logo[7][20] = 9'b111101101;
assign reset_logo[7][21] = 9'b111101101;
assign reset_logo[7][22] = 9'b111101101;
assign reset_logo[7][23] = 9'b111101001;
assign reset_logo[7][24] = 9'b111101101;
assign reset_logo[7][25] = 9'b111101101;
assign reset_logo[7][26] = 9'b111101001;
assign reset_logo[7][27] = 9'b111101001;
assign reset_logo[7][28] = 9'b101101101;
assign reset_logo[7][29] = 9'b101001001;
assign reset_logo[7][30] = 9'b101001001;
assign reset_logo[7][31] = 9'b101001001;
assign reset_logo[7][32] = 9'b101101101;
assign reset_logo[7][33] = 9'b101001001;
assign reset_logo[7][34] = 9'b101001001;
assign reset_logo[7][35] = 9'b101001001;
assign reset_logo[8][3] = 9'b100100100;
assign reset_logo[8][4] = 9'b100100100;
assign reset_logo[8][5] = 9'b100100100;
assign reset_logo[8][6] = 9'b101001001;
assign reset_logo[8][7] = 9'b101001001;
assign reset_logo[8][8] = 9'b101101001;
assign reset_logo[8][9] = 9'b101101101;
assign reset_logo[8][10] = 9'b110010001;
assign reset_logo[8][11] = 9'b111101001;
assign reset_logo[8][12] = 9'b111100100;
assign reset_logo[8][13] = 9'b111100100;
assign reset_logo[8][14] = 9'b111101000;
assign reset_logo[8][15] = 9'b111101101;
assign reset_logo[8][16] = 9'b111110001;
assign reset_logo[8][17] = 9'b111111110;
assign reset_logo[8][18] = 9'b111111111;
assign reset_logo[8][19] = 9'b111111111;
assign reset_logo[8][20] = 9'b111111111;
assign reset_logo[8][21] = 9'b111111111;
assign reset_logo[8][22] = 9'b111111111;
assign reset_logo[8][23] = 9'b111111110;
assign reset_logo[8][24] = 9'b111110001;
assign reset_logo[8][25] = 9'b111101101;
assign reset_logo[8][26] = 9'b111101101;
assign reset_logo[8][27] = 9'b111101101;
assign reset_logo[8][28] = 9'b111101001;
assign reset_logo[8][29] = 9'b110001001;
assign reset_logo[8][30] = 9'b101001001;
assign reset_logo[8][31] = 9'b101001001;
assign reset_logo[8][32] = 9'b101001001;
assign reset_logo[8][33] = 9'b101101101;
assign reset_logo[8][34] = 9'b101001001;
assign reset_logo[8][35] = 9'b101001001;
assign reset_logo[8][36] = 9'b100100100;
assign reset_logo[9][3] = 9'b100100100;
assign reset_logo[9][4] = 9'b100100100;
assign reset_logo[9][5] = 9'b101001001;
assign reset_logo[9][6] = 9'b101001001;
assign reset_logo[9][7] = 9'b101101001;
assign reset_logo[9][8] = 9'b101101101;
assign reset_logo[9][9] = 9'b110010001;
assign reset_logo[9][10] = 9'b111101000;
assign reset_logo[9][11] = 9'b111100100;
assign reset_logo[9][12] = 9'b111100100;
assign reset_logo[9][13] = 9'b111101101;
assign reset_logo[9][14] = 9'b111110101;
assign reset_logo[9][15] = 9'b111111110;
assign reset_logo[9][16] = 9'b111110110;
assign reset_logo[9][17] = 9'b111110001;
assign reset_logo[9][18] = 9'b111110001;
assign reset_logo[9][19] = 9'b111110001;
assign reset_logo[9][20] = 9'b111110001;
assign reset_logo[9][21] = 9'b111110110;
assign reset_logo[9][22] = 9'b111110110;
assign reset_logo[9][23] = 9'b111111111;
assign reset_logo[9][24] = 9'b111111111;
assign reset_logo[9][25] = 9'b111111111;
assign reset_logo[9][26] = 9'b111110001;
assign reset_logo[9][27] = 9'b111101101;
assign reset_logo[9][28] = 9'b111101101;
assign reset_logo[9][29] = 9'b111101001;
assign reset_logo[9][30] = 9'b110001001;
assign reset_logo[9][31] = 9'b101001001;
assign reset_logo[9][32] = 9'b101001000;
assign reset_logo[9][33] = 9'b101001001;
assign reset_logo[9][34] = 9'b101001001;
assign reset_logo[9][35] = 9'b101001001;
assign reset_logo[9][36] = 9'b101001001;
assign reset_logo[10][2] = 9'b100100100;
assign reset_logo[10][3] = 9'b100100100;
assign reset_logo[10][4] = 9'b101001001;
assign reset_logo[10][5] = 9'b101001001;
assign reset_logo[10][6] = 9'b101101001;
assign reset_logo[10][7] = 9'b101101101;
assign reset_logo[10][8] = 9'b110010001;
assign reset_logo[10][9] = 9'b111101000;
assign reset_logo[10][10] = 9'b111100100;
assign reset_logo[10][11] = 9'b111100100;
assign reset_logo[10][12] = 9'b111101000;
assign reset_logo[10][13] = 9'b111101101;
assign reset_logo[10][14] = 9'b111101101;
assign reset_logo[10][15] = 9'b111101000;
assign reset_logo[10][16] = 9'b111101000;
assign reset_logo[10][17] = 9'b111101000;
assign reset_logo[10][18] = 9'b111101001;
assign reset_logo[10][19] = 9'b111101101;
assign reset_logo[10][20] = 9'b111101101;
assign reset_logo[10][21] = 9'b111101101;
assign reset_logo[10][22] = 9'b111101101;
assign reset_logo[10][23] = 9'b111101101;
assign reset_logo[10][24] = 9'b111101101;
assign reset_logo[10][25] = 9'b111110001;
assign reset_logo[10][26] = 9'b111110110;
assign reset_logo[10][27] = 9'b111110001;
assign reset_logo[10][28] = 9'b111101101;
assign reset_logo[10][29] = 9'b111101101;
assign reset_logo[10][30] = 9'b111101001;
assign reset_logo[10][31] = 9'b101101001;
assign reset_logo[10][32] = 9'b101001000;
assign reset_logo[10][33] = 9'b101001000;
assign reset_logo[10][34] = 9'b101001001;
assign reset_logo[10][35] = 9'b101001001;
assign reset_logo[10][36] = 9'b101001000;
assign reset_logo[10][37] = 9'b100100100;
assign reset_logo[11][2] = 9'b100100100;
assign reset_logo[11][3] = 9'b101001000;
assign reset_logo[11][4] = 9'b101001001;
assign reset_logo[11][5] = 9'b101001001;
assign reset_logo[11][6] = 9'b101101101;
assign reset_logo[11][7] = 9'b101110001;
assign reset_logo[11][8] = 9'b111101001;
assign reset_logo[11][9] = 9'b111100100;
assign reset_logo[11][10] = 9'b111100100;
assign reset_logo[11][11] = 9'b111100100;
assign reset_logo[11][12] = 9'b111101000;
assign reset_logo[11][13] = 9'b111101000;
assign reset_logo[11][14] = 9'b111101000;
assign reset_logo[11][15] = 9'b111101000;
assign reset_logo[11][16] = 9'b111101001;
assign reset_logo[11][17] = 9'b111101001;
assign reset_logo[11][18] = 9'b111101101;
assign reset_logo[11][19] = 9'b111101101;
assign reset_logo[11][20] = 9'b111101101;
assign reset_logo[11][21] = 9'b111101101;
assign reset_logo[11][22] = 9'b111101101;
assign reset_logo[11][23] = 9'b111101101;
assign reset_logo[11][24] = 9'b111110001;
assign reset_logo[11][25] = 9'b111101101;
assign reset_logo[11][26] = 9'b111101101;
assign reset_logo[11][27] = 9'b111101101;
assign reset_logo[11][28] = 9'b111101101;
assign reset_logo[11][29] = 9'b111101101;
assign reset_logo[11][30] = 9'b111101101;
assign reset_logo[11][31] = 9'b111101001;
assign reset_logo[11][32] = 9'b101101001;
assign reset_logo[11][33] = 9'b101001000;
assign reset_logo[11][34] = 9'b101001000;
assign reset_logo[11][35] = 9'b101001000;
assign reset_logo[11][36] = 9'b100100100;
assign reset_logo[11][37] = 9'b101001000;
assign reset_logo[12][1] = 9'b100100100;
assign reset_logo[12][2] = 9'b101001000;
assign reset_logo[12][3] = 9'b101001001;
assign reset_logo[12][4] = 9'b101001001;
assign reset_logo[12][5] = 9'b101101101;
assign reset_logo[12][6] = 9'b101101101;
assign reset_logo[12][7] = 9'b110101101;
assign reset_logo[12][8] = 9'b111100100;
assign reset_logo[12][9] = 9'b111100100;
assign reset_logo[12][10] = 9'b111100100;
assign reset_logo[12][11] = 9'b111100100;
assign reset_logo[12][12] = 9'b111101000;
assign reset_logo[12][13] = 9'b111101000;
assign reset_logo[12][14] = 9'b111101000;
assign reset_logo[12][15] = 9'b111101000;
assign reset_logo[12][16] = 9'b111101001;
assign reset_logo[12][17] = 9'b111101101;
assign reset_logo[12][18] = 9'b111101101;
assign reset_logo[12][19] = 9'b111101101;
assign reset_logo[12][20] = 9'b111101101;
assign reset_logo[12][21] = 9'b111101101;
assign reset_logo[12][22] = 9'b111110001;
assign reset_logo[12][23] = 9'b111110001;
assign reset_logo[12][24] = 9'b111110001;
assign reset_logo[12][25] = 9'b111110001;
assign reset_logo[12][26] = 9'b111110001;
assign reset_logo[12][27] = 9'b111101101;
assign reset_logo[12][28] = 9'b111101101;
assign reset_logo[12][29] = 9'b111101101;
assign reset_logo[12][30] = 9'b111101101;
assign reset_logo[12][31] = 9'b111101101;
assign reset_logo[12][32] = 9'b110101001;
assign reset_logo[12][33] = 9'b101001000;
assign reset_logo[12][34] = 9'b100100100;
assign reset_logo[12][35] = 9'b100100100;
assign reset_logo[12][36] = 9'b100100100;
assign reset_logo[12][37] = 9'b100100100;
assign reset_logo[12][38] = 9'b100100100;
assign reset_logo[13][1] = 9'b101001000;
assign reset_logo[13][2] = 9'b101001000;
assign reset_logo[13][3] = 9'b101001001;
assign reset_logo[13][4] = 9'b101101101;
assign reset_logo[13][5] = 9'b101101101;
assign reset_logo[13][6] = 9'b110010001;
assign reset_logo[13][7] = 9'b111101000;
assign reset_logo[13][8] = 9'b111100000;
assign reset_logo[13][9] = 9'b111100100;
assign reset_logo[13][10] = 9'b111100100;
assign reset_logo[13][11] = 9'b111100100;
assign reset_logo[13][12] = 9'b111101000;
assign reset_logo[13][13] = 9'b111101000;
assign reset_logo[13][14] = 9'b111101000;
assign reset_logo[13][15] = 9'b111101000;
assign reset_logo[13][16] = 9'b111101001;
assign reset_logo[13][17] = 9'b111101101;
assign reset_logo[13][18] = 9'b111101101;
assign reset_logo[13][19] = 9'b111101101;
assign reset_logo[13][20] = 9'b111101101;
assign reset_logo[13][21] = 9'b111101101;
assign reset_logo[13][22] = 9'b111110001;
assign reset_logo[13][23] = 9'b111110001;
assign reset_logo[13][24] = 9'b111110001;
assign reset_logo[13][25] = 9'b111110001;
assign reset_logo[13][26] = 9'b111110001;
assign reset_logo[13][27] = 9'b111110001;
assign reset_logo[13][28] = 9'b111101101;
assign reset_logo[13][29] = 9'b111101101;
assign reset_logo[13][30] = 9'b111101101;
assign reset_logo[13][31] = 9'b111101101;
assign reset_logo[13][32] = 9'b111101001;
assign reset_logo[13][33] = 9'b101101000;
assign reset_logo[13][34] = 9'b100100100;
assign reset_logo[13][35] = 9'b100100100;
assign reset_logo[13][36] = 9'b100100100;
assign reset_logo[13][37] = 9'b100100100;
assign reset_logo[13][38] = 9'b100100100;
assign reset_logo[14][1] = 9'b101001000;
assign reset_logo[14][2] = 9'b101001001;
assign reset_logo[14][3] = 9'b101101101;
assign reset_logo[14][4] = 9'b101101101;
assign reset_logo[14][5] = 9'b101101101;
assign reset_logo[14][6] = 9'b110101101;
assign reset_logo[14][7] = 9'b111100100;
assign reset_logo[14][8] = 9'b111100100;
assign reset_logo[14][9] = 9'b111100100;
assign reset_logo[14][10] = 9'b111100100;
assign reset_logo[14][11] = 9'b111100100;
assign reset_logo[14][12] = 9'b111101000;
assign reset_logo[14][13] = 9'b111101000;
assign reset_logo[14][14] = 9'b111101000;
assign reset_logo[14][15] = 9'b111101000;
assign reset_logo[14][16] = 9'b111101001;
assign reset_logo[14][17] = 9'b111101101;
assign reset_logo[14][18] = 9'b111101101;
assign reset_logo[14][19] = 9'b111101101;
assign reset_logo[14][20] = 9'b111101101;
assign reset_logo[14][21] = 9'b111101101;
assign reset_logo[14][22] = 9'b111110001;
assign reset_logo[14][23] = 9'b111110001;
assign reset_logo[14][24] = 9'b111110001;
assign reset_logo[14][25] = 9'b111110001;
assign reset_logo[14][26] = 9'b111110001;
assign reset_logo[14][27] = 9'b111110001;
assign reset_logo[14][28] = 9'b111101101;
assign reset_logo[14][29] = 9'b111101101;
assign reset_logo[14][30] = 9'b111101101;
assign reset_logo[14][31] = 9'b111101101;
assign reset_logo[14][32] = 9'b111101001;
assign reset_logo[14][33] = 9'b110101001;
assign reset_logo[14][34] = 9'b100100100;
assign reset_logo[14][35] = 9'b100100100;
assign reset_logo[14][36] = 9'b100100100;
assign reset_logo[14][37] = 9'b100100100;
assign reset_logo[14][38] = 9'b100100100;
assign reset_logo[15][0] = 9'b101001000;
assign reset_logo[15][1] = 9'b101001001;
assign reset_logo[15][2] = 9'b101001001;
assign reset_logo[15][3] = 9'b101101101;
assign reset_logo[15][4] = 9'b101101101;
assign reset_logo[15][5] = 9'b110010001;
assign reset_logo[15][6] = 9'b111101101;
assign reset_logo[15][7] = 9'b111100000;
assign reset_logo[15][8] = 9'b111100100;
assign reset_logo[15][9] = 9'b111100100;
assign reset_logo[15][10] = 9'b111100100;
assign reset_logo[15][11] = 9'b111100100;
assign reset_logo[15][12] = 9'b111101000;
assign reset_logo[15][13] = 9'b111101000;
assign reset_logo[15][14] = 9'b111101000;
assign reset_logo[15][15] = 9'b111101000;
assign reset_logo[15][16] = 9'b111101000;
assign reset_logo[15][17] = 9'b111101101;
assign reset_logo[15][18] = 9'b111101101;
assign reset_logo[15][19] = 9'b111101101;
assign reset_logo[15][20] = 9'b111101101;
assign reset_logo[15][21] = 9'b111101101;
assign reset_logo[15][22] = 9'b111110001;
assign reset_logo[15][23] = 9'b111110001;
assign reset_logo[15][24] = 9'b111110001;
assign reset_logo[15][25] = 9'b111110001;
assign reset_logo[15][26] = 9'b111110001;
assign reset_logo[15][27] = 9'b111101101;
assign reset_logo[15][28] = 9'b111101101;
assign reset_logo[15][29] = 9'b111101101;
assign reset_logo[15][30] = 9'b111101101;
assign reset_logo[15][31] = 9'b111101101;
assign reset_logo[15][32] = 9'b111101101;
assign reset_logo[15][33] = 9'b111101001;
assign reset_logo[15][34] = 9'b101001000;
assign reset_logo[15][35] = 9'b100100000;
assign reset_logo[15][36] = 9'b100100000;
assign reset_logo[15][37] = 9'b100100100;
assign reset_logo[15][38] = 9'b100100100;
assign reset_logo[15][39] = 9'b100000000;
assign reset_logo[16][0] = 9'b101001000;
assign reset_logo[16][1] = 9'b101001001;
assign reset_logo[16][2] = 9'b101101101;
assign reset_logo[16][3] = 9'b101101101;
assign reset_logo[16][4] = 9'b101101101;
assign reset_logo[16][5] = 9'b110010001;
assign reset_logo[16][6] = 9'b111101000;
assign reset_logo[16][7] = 9'b111100000;
assign reset_logo[16][8] = 9'b111100100;
assign reset_logo[16][9] = 9'b111101000;
assign reset_logo[16][10] = 9'b111101001;
assign reset_logo[16][11] = 9'b111101000;
assign reset_logo[16][12] = 9'b111100100;
assign reset_logo[16][13] = 9'b111101000;
assign reset_logo[16][14] = 9'b111101101;
assign reset_logo[16][15] = 9'b111101101;
assign reset_logo[16][16] = 9'b111101101;
assign reset_logo[16][17] = 9'b111101101;
assign reset_logo[16][18] = 9'b111101101;
assign reset_logo[16][19] = 9'b111110001;
assign reset_logo[16][20] = 9'b111110001;
assign reset_logo[16][21] = 9'b111110001;
assign reset_logo[16][22] = 9'b111110001;
assign reset_logo[16][23] = 9'b111110001;
assign reset_logo[16][24] = 9'b111110001;
assign reset_logo[16][25] = 9'b111110001;
assign reset_logo[16][26] = 9'b111110001;
assign reset_logo[16][27] = 9'b111110001;
assign reset_logo[16][28] = 9'b111110001;
assign reset_logo[16][29] = 9'b111110001;
assign reset_logo[16][30] = 9'b111110001;
assign reset_logo[16][31] = 9'b111101101;
assign reset_logo[16][32] = 9'b111101001;
assign reset_logo[16][33] = 9'b111101001;
assign reset_logo[16][34] = 9'b101101000;
assign reset_logo[16][35] = 9'b100100100;
assign reset_logo[16][36] = 9'b100000000;
assign reset_logo[16][37] = 9'b100000000;
assign reset_logo[16][38] = 9'b100000000;
assign reset_logo[16][39] = 9'b100000000;
assign reset_logo[17][0] = 9'b101001001;
assign reset_logo[17][1] = 9'b101001001;
assign reset_logo[17][2] = 9'b101101101;
assign reset_logo[17][3] = 9'b101101101;
assign reset_logo[17][4] = 9'b101101101;
assign reset_logo[17][5] = 9'b110010001;
assign reset_logo[17][6] = 9'b111100100;
assign reset_logo[17][7] = 9'b111100000;
assign reset_logo[17][8] = 9'b111101101;
assign reset_logo[17][9] = 9'b111111111;
assign reset_logo[17][10] = 9'b111111110;
assign reset_logo[17][11] = 9'b111111111;
assign reset_logo[17][12] = 9'b111101101;
assign reset_logo[17][13] = 9'b111101101;
assign reset_logo[17][14] = 9'b111111111;
assign reset_logo[17][15] = 9'b111111111;
assign reset_logo[17][16] = 9'b111111111;
assign reset_logo[17][17] = 9'b111101101;
assign reset_logo[17][18] = 9'b111110110;
assign reset_logo[17][19] = 9'b111111111;
assign reset_logo[17][20] = 9'b111111111;
assign reset_logo[17][21] = 9'b111110110;
assign reset_logo[17][22] = 9'b111110001;
assign reset_logo[17][23] = 9'b111111111;
assign reset_logo[17][24] = 9'b111111111;
assign reset_logo[17][25] = 9'b111111111;
assign reset_logo[17][26] = 9'b111110110;
assign reset_logo[17][27] = 9'b111111111;
assign reset_logo[17][28] = 9'b111111111;
assign reset_logo[17][29] = 9'b111111111;
assign reset_logo[17][30] = 9'b111111111;
assign reset_logo[17][31] = 9'b111110001;
assign reset_logo[17][32] = 9'b111101000;
assign reset_logo[17][33] = 9'b111101000;
assign reset_logo[17][34] = 9'b110001001;
assign reset_logo[17][35] = 9'b100100100;
assign reset_logo[17][36] = 9'b100000000;
assign reset_logo[17][37] = 9'b100000000;
assign reset_logo[17][38] = 9'b100000000;
assign reset_logo[17][39] = 9'b100000000;
assign reset_logo[18][0] = 9'b101001001;
assign reset_logo[18][1] = 9'b101001001;
assign reset_logo[18][2] = 9'b101101101;
assign reset_logo[18][3] = 9'b101101101;
assign reset_logo[18][4] = 9'b110010001;
assign reset_logo[18][5] = 9'b110010001;
assign reset_logo[18][6] = 9'b111100100;
assign reset_logo[18][7] = 9'b111100000;
assign reset_logo[18][8] = 9'b111101101;
assign reset_logo[18][9] = 9'b111111111;
assign reset_logo[18][10] = 9'b111100000;
assign reset_logo[18][11] = 9'b111111111;
assign reset_logo[18][12] = 9'b111111111;
assign reset_logo[18][13] = 9'b111101001;
assign reset_logo[18][14] = 9'b111111111;
assign reset_logo[18][15] = 9'b111101001;
assign reset_logo[18][16] = 9'b111101000;
assign reset_logo[18][17] = 9'b111101101;
assign reset_logo[18][18] = 9'b111111111;
assign reset_logo[18][19] = 9'b111110110;
assign reset_logo[18][20] = 9'b111101000;
assign reset_logo[18][21] = 9'b111101101;
assign reset_logo[18][22] = 9'b111101101;
assign reset_logo[18][23] = 9'b111111111;
assign reset_logo[18][24] = 9'b111110001;
assign reset_logo[18][25] = 9'b111101101;
assign reset_logo[18][26] = 9'b111101101;
assign reset_logo[18][27] = 9'b111101101;
assign reset_logo[18][28] = 9'b111110110;
assign reset_logo[18][29] = 9'b111111111;
assign reset_logo[18][30] = 9'b111101101;
assign reset_logo[18][31] = 9'b111101001;
assign reset_logo[18][32] = 9'b111101001;
assign reset_logo[18][33] = 9'b111101000;
assign reset_logo[18][34] = 9'b110001001;
assign reset_logo[18][35] = 9'b100100100;
assign reset_logo[18][36] = 9'b100100000;
assign reset_logo[18][37] = 9'b100000000;
assign reset_logo[18][38] = 9'b100000000;
assign reset_logo[18][39] = 9'b100000000;
assign reset_logo[19][0] = 9'b101001001;
assign reset_logo[19][1] = 9'b101101101;
assign reset_logo[19][2] = 9'b101101101;
assign reset_logo[19][3] = 9'b110010001;
assign reset_logo[19][4] = 9'b110010001;
assign reset_logo[19][5] = 9'b110110001;
assign reset_logo[19][6] = 9'b111100100;
assign reset_logo[19][7] = 9'b111100000;
assign reset_logo[19][8] = 9'b111101101;
assign reset_logo[19][9] = 9'b111111111;
assign reset_logo[19][10] = 9'b111110110;
assign reset_logo[19][11] = 9'b111111111;
assign reset_logo[19][12] = 9'b111101101;
assign reset_logo[19][13] = 9'b111101001;
assign reset_logo[19][14] = 9'b111111111;
assign reset_logo[19][15] = 9'b111111111;
assign reset_logo[19][16] = 9'b111111111;
assign reset_logo[19][17] = 9'b111101101;
assign reset_logo[19][18] = 9'b111110001;
assign reset_logo[19][19] = 9'b111111111;
assign reset_logo[19][20] = 9'b111110110;
assign reset_logo[19][21] = 9'b111101101;
assign reset_logo[19][22] = 9'b111101101;
assign reset_logo[19][23] = 9'b111111111;
assign reset_logo[19][24] = 9'b111111111;
assign reset_logo[19][25] = 9'b111111111;
assign reset_logo[19][26] = 9'b111110001;
assign reset_logo[19][27] = 9'b111101001;
assign reset_logo[19][28] = 9'b111110110;
assign reset_logo[19][29] = 9'b111111111;
assign reset_logo[19][30] = 9'b111101101;
assign reset_logo[19][31] = 9'b111101001;
assign reset_logo[19][32] = 9'b111101000;
assign reset_logo[19][33] = 9'b111101000;
assign reset_logo[19][34] = 9'b110001001;
assign reset_logo[19][35] = 9'b100100100;
assign reset_logo[19][36] = 9'b100100100;
assign reset_logo[19][37] = 9'b100000000;
assign reset_logo[19][38] = 9'b100000000;
assign reset_logo[19][39] = 9'b100000000;
assign reset_logo[20][0] = 9'b101001001;
assign reset_logo[20][1] = 9'b101001001;
assign reset_logo[20][2] = 9'b101101101;
assign reset_logo[20][3] = 9'b110010001;
assign reset_logo[20][4] = 9'b110010001;
assign reset_logo[20][5] = 9'b110010001;
assign reset_logo[20][6] = 9'b111100100;
assign reset_logo[20][7] = 9'b111100000;
assign reset_logo[20][8] = 9'b111101101;
assign reset_logo[20][9] = 9'b111111111;
assign reset_logo[20][10] = 9'b111111111;
assign reset_logo[20][11] = 9'b111110010;
assign reset_logo[20][12] = 9'b111100000;
assign reset_logo[20][13] = 9'b111101101;
assign reset_logo[20][14] = 9'b111111111;
assign reset_logo[20][15] = 9'b111101101;
assign reset_logo[20][16] = 9'b111101101;
assign reset_logo[20][17] = 9'b111101001;
assign reset_logo[20][18] = 9'b111101000;
assign reset_logo[20][19] = 9'b111101101;
assign reset_logo[20][20] = 9'b111111111;
assign reset_logo[20][21] = 9'b111111111;
assign reset_logo[20][22] = 9'b111101101;
assign reset_logo[20][23] = 9'b111111111;
assign reset_logo[20][24] = 9'b111110010;
assign reset_logo[20][25] = 9'b111101101;
assign reset_logo[20][26] = 9'b111101101;
assign reset_logo[20][27] = 9'b111101001;
assign reset_logo[20][28] = 9'b111110010;
assign reset_logo[20][29] = 9'b111111111;
assign reset_logo[20][30] = 9'b111101001;
assign reset_logo[20][31] = 9'b111101000;
assign reset_logo[20][32] = 9'b111101000;
assign reset_logo[20][33] = 9'b111101000;
assign reset_logo[20][34] = 9'b110001001;
assign reset_logo[20][35] = 9'b100101000;
assign reset_logo[20][36] = 9'b100100100;
assign reset_logo[20][37] = 9'b100000000;
assign reset_logo[20][38] = 9'b100000000;
assign reset_logo[20][39] = 9'b100000000;
assign reset_logo[21][0] = 9'b101001001;
assign reset_logo[21][1] = 9'b101001001;
assign reset_logo[21][2] = 9'b101101101;
assign reset_logo[21][3] = 9'b101101101;
assign reset_logo[21][4] = 9'b101101101;
assign reset_logo[21][5] = 9'b110010001;
assign reset_logo[21][6] = 9'b111100100;
assign reset_logo[21][7] = 9'b111100000;
assign reset_logo[21][8] = 9'b111101101;
assign reset_logo[21][9] = 9'b111111111;
assign reset_logo[21][10] = 9'b111101000;
assign reset_logo[21][11] = 9'b111111111;
assign reset_logo[21][12] = 9'b111101101;
assign reset_logo[21][13] = 9'b111101001;
assign reset_logo[21][14] = 9'b111111111;
assign reset_logo[21][15] = 9'b111101101;
assign reset_logo[21][16] = 9'b111101001;
assign reset_logo[21][17] = 9'b111101001;
assign reset_logo[21][18] = 9'b111101101;
assign reset_logo[21][19] = 9'b111101101;
assign reset_logo[21][20] = 9'b111110010;
assign reset_logo[21][21] = 9'b111111111;
assign reset_logo[21][22] = 9'b111101101;
assign reset_logo[21][23] = 9'b111111111;
assign reset_logo[21][24] = 9'b111110001;
assign reset_logo[21][25] = 9'b111101101;
assign reset_logo[21][26] = 9'b111101101;
assign reset_logo[21][27] = 9'b111101000;
assign reset_logo[21][28] = 9'b111110110;
assign reset_logo[21][29] = 9'b111111111;
assign reset_logo[21][30] = 9'b111101001;
assign reset_logo[21][31] = 9'b111101000;
assign reset_logo[21][32] = 9'b111101000;
assign reset_logo[21][33] = 9'b111101000;
assign reset_logo[21][34] = 9'b110001001;
assign reset_logo[21][35] = 9'b100101000;
assign reset_logo[21][36] = 9'b100100100;
assign reset_logo[21][37] = 9'b100100100;
assign reset_logo[21][38] = 9'b100000000;
assign reset_logo[21][39] = 9'b100000000;
assign reset_logo[22][0] = 9'b101001001;
assign reset_logo[22][1] = 9'b101001001;
assign reset_logo[22][2] = 9'b101101101;
assign reset_logo[22][3] = 9'b101101101;
assign reset_logo[22][4] = 9'b101101101;
assign reset_logo[22][5] = 9'b110010001;
assign reset_logo[22][6] = 9'b111101000;
assign reset_logo[22][7] = 9'b111100000;
assign reset_logo[22][8] = 9'b111101001;
assign reset_logo[22][9] = 9'b111111110;
assign reset_logo[22][10] = 9'b111100000;
assign reset_logo[22][11] = 9'b111101101;
assign reset_logo[22][12] = 9'b111110110;
assign reset_logo[22][13] = 9'b111101001;
assign reset_logo[22][14] = 9'b111111111;
assign reset_logo[22][15] = 9'b111111111;
assign reset_logo[22][16] = 9'b111111111;
assign reset_logo[22][17] = 9'b111101101;
assign reset_logo[22][18] = 9'b111110001;
assign reset_logo[22][19] = 9'b111111111;
assign reset_logo[22][20] = 9'b111111111;
assign reset_logo[22][21] = 9'b111110001;
assign reset_logo[22][22] = 9'b111101001;
assign reset_logo[22][23] = 9'b111111111;
assign reset_logo[22][24] = 9'b111111111;
assign reset_logo[22][25] = 9'b111111111;
assign reset_logo[22][26] = 9'b111110001;
assign reset_logo[22][27] = 9'b111101000;
assign reset_logo[22][28] = 9'b111110001;
assign reset_logo[22][29] = 9'b111111111;
assign reset_logo[22][30] = 9'b111101000;
assign reset_logo[22][31] = 9'b111101000;
assign reset_logo[22][32] = 9'b111101000;
assign reset_logo[22][33] = 9'b111101000;
assign reset_logo[22][34] = 9'b110001001;
assign reset_logo[22][35] = 9'b101001000;
assign reset_logo[22][36] = 9'b100100100;
assign reset_logo[22][37] = 9'b100100100;
assign reset_logo[22][38] = 9'b100000000;
assign reset_logo[22][39] = 9'b100000000;
assign reset_logo[23][0] = 9'b101101101;
assign reset_logo[23][1] = 9'b101101101;
assign reset_logo[23][2] = 9'b101101101;
assign reset_logo[23][3] = 9'b101001001;
assign reset_logo[23][4] = 9'b101101101;
assign reset_logo[23][5] = 9'b101110001;
assign reset_logo[23][6] = 9'b111101001;
assign reset_logo[23][7] = 9'b111100000;
assign reset_logo[23][8] = 9'b111100000;
assign reset_logo[23][9] = 9'b111100000;
assign reset_logo[23][10] = 9'b111100100;
assign reset_logo[23][11] = 9'b111100000;
assign reset_logo[23][12] = 9'b111100100;
assign reset_logo[23][13] = 9'b111100100;
assign reset_logo[23][14] = 9'b111100100;
assign reset_logo[23][15] = 9'b111100100;
assign reset_logo[23][16] = 9'b111101000;
assign reset_logo[23][17] = 9'b111101000;
assign reset_logo[23][18] = 9'b111101000;
assign reset_logo[23][19] = 9'b111101000;
assign reset_logo[23][20] = 9'b111101000;
assign reset_logo[23][21] = 9'b111101000;
assign reset_logo[23][22] = 9'b111101000;
assign reset_logo[23][23] = 9'b111101000;
assign reset_logo[23][24] = 9'b111101000;
assign reset_logo[23][25] = 9'b111101000;
assign reset_logo[23][26] = 9'b111101000;
assign reset_logo[23][27] = 9'b111101000;
assign reset_logo[23][28] = 9'b111101000;
assign reset_logo[23][29] = 9'b111101000;
assign reset_logo[23][30] = 9'b111101000;
assign reset_logo[23][31] = 9'b111101000;
assign reset_logo[23][32] = 9'b111101000;
assign reset_logo[23][33] = 9'b111101000;
assign reset_logo[23][34] = 9'b101101001;
assign reset_logo[23][35] = 9'b101001000;
assign reset_logo[23][36] = 9'b100100100;
assign reset_logo[23][37] = 9'b100100100;
assign reset_logo[23][38] = 9'b100000000;
assign reset_logo[23][39] = 9'b100000000;
assign reset_logo[24][0] = 9'b101101101;
assign reset_logo[24][1] = 9'b101101101;
assign reset_logo[24][2] = 9'b101101101;
assign reset_logo[24][3] = 9'b101101101;
assign reset_logo[24][4] = 9'b101001001;
assign reset_logo[24][5] = 9'b101101101;
assign reset_logo[24][6] = 9'b111101101;
assign reset_logo[24][7] = 9'b111100000;
assign reset_logo[24][8] = 9'b111100000;
assign reset_logo[24][9] = 9'b111100000;
assign reset_logo[24][10] = 9'b111100100;
assign reset_logo[24][11] = 9'b111100100;
assign reset_logo[24][12] = 9'b111100100;
assign reset_logo[24][13] = 9'b111100100;
assign reset_logo[24][14] = 9'b111100100;
assign reset_logo[24][15] = 9'b111100100;
assign reset_logo[24][16] = 9'b111100100;
assign reset_logo[24][17] = 9'b111101000;
assign reset_logo[24][18] = 9'b111101000;
assign reset_logo[24][19] = 9'b111101000;
assign reset_logo[24][20] = 9'b111101000;
assign reset_logo[24][21] = 9'b111101000;
assign reset_logo[24][22] = 9'b111101000;
assign reset_logo[24][23] = 9'b111101000;
assign reset_logo[24][24] = 9'b111101000;
assign reset_logo[24][25] = 9'b111101000;
assign reset_logo[24][26] = 9'b111101000;
assign reset_logo[24][27] = 9'b111101000;
assign reset_logo[24][28] = 9'b111101000;
assign reset_logo[24][29] = 9'b111101000;
assign reset_logo[24][30] = 9'b111101000;
assign reset_logo[24][31] = 9'b111101000;
assign reset_logo[24][32] = 9'b111100100;
assign reset_logo[24][33] = 9'b111101001;
assign reset_logo[24][34] = 9'b101001001;
assign reset_logo[24][35] = 9'b101001000;
assign reset_logo[24][36] = 9'b100100100;
assign reset_logo[24][37] = 9'b100100100;
assign reset_logo[24][38] = 9'b100000000;
assign reset_logo[24][39] = 9'b100000000;
assign reset_logo[25][1] = 9'b101101101;
assign reset_logo[25][2] = 9'b101101101;
assign reset_logo[25][3] = 9'b101101101;
assign reset_logo[25][4] = 9'b101101001;
assign reset_logo[25][5] = 9'b101001001;
assign reset_logo[25][6] = 9'b110010001;
assign reset_logo[25][7] = 9'b111101000;
assign reset_logo[25][8] = 9'b111100000;
assign reset_logo[25][9] = 9'b111100100;
assign reset_logo[25][10] = 9'b111100100;
assign reset_logo[25][11] = 9'b111100100;
assign reset_logo[25][12] = 9'b111100100;
assign reset_logo[25][13] = 9'b111100100;
assign reset_logo[25][14] = 9'b111100100;
assign reset_logo[25][15] = 9'b111100100;
assign reset_logo[25][16] = 9'b111100100;
assign reset_logo[25][17] = 9'b111100100;
assign reset_logo[25][18] = 9'b111100100;
assign reset_logo[25][19] = 9'b111101000;
assign reset_logo[25][20] = 9'b111101000;
assign reset_logo[25][21] = 9'b111101000;
assign reset_logo[25][22] = 9'b111101000;
assign reset_logo[25][23] = 9'b111101000;
assign reset_logo[25][24] = 9'b111101000;
assign reset_logo[25][25] = 9'b111101000;
assign reset_logo[25][26] = 9'b111101000;
assign reset_logo[25][27] = 9'b111101000;
assign reset_logo[25][28] = 9'b111101000;
assign reset_logo[25][29] = 9'b111101000;
assign reset_logo[25][30] = 9'b111101000;
assign reset_logo[25][31] = 9'b111100100;
assign reset_logo[25][32] = 9'b111100100;
assign reset_logo[25][33] = 9'b110001101;
assign reset_logo[25][34] = 9'b101001001;
assign reset_logo[25][35] = 9'b101001001;
assign reset_logo[25][36] = 9'b101001000;
assign reset_logo[25][37] = 9'b100100100;
assign reset_logo[25][38] = 9'b100000000;
assign reset_logo[26][1] = 9'b101101101;
assign reset_logo[26][2] = 9'b101101101;
assign reset_logo[26][3] = 9'b101101101;
assign reset_logo[26][4] = 9'b101101101;
assign reset_logo[26][5] = 9'b101001001;
assign reset_logo[26][6] = 9'b101101101;
assign reset_logo[26][7] = 9'b111101101;
assign reset_logo[26][8] = 9'b111100000;
assign reset_logo[26][9] = 9'b111100000;
assign reset_logo[26][10] = 9'b111100100;
assign reset_logo[26][11] = 9'b111100100;
assign reset_logo[26][12] = 9'b111100100;
assign reset_logo[26][13] = 9'b111100100;
assign reset_logo[26][14] = 9'b111100100;
assign reset_logo[26][15] = 9'b111100100;
assign reset_logo[26][16] = 9'b111100100;
assign reset_logo[26][17] = 9'b111100100;
assign reset_logo[26][18] = 9'b111100100;
assign reset_logo[26][19] = 9'b111100100;
assign reset_logo[26][20] = 9'b111100100;
assign reset_logo[26][21] = 9'b111101000;
assign reset_logo[26][22] = 9'b111101000;
assign reset_logo[26][23] = 9'b111101000;
assign reset_logo[26][24] = 9'b111101000;
assign reset_logo[26][25] = 9'b111101000;
assign reset_logo[26][26] = 9'b111101000;
assign reset_logo[26][27] = 9'b111101000;
assign reset_logo[26][28] = 9'b111100100;
assign reset_logo[26][29] = 9'b111100100;
assign reset_logo[26][30] = 9'b111100100;
assign reset_logo[26][31] = 9'b111100100;
assign reset_logo[26][32] = 9'b111101001;
assign reset_logo[26][33] = 9'b101101101;
assign reset_logo[26][34] = 9'b101101101;
assign reset_logo[26][35] = 9'b101001001;
assign reset_logo[26][36] = 9'b101001001;
assign reset_logo[26][37] = 9'b100100100;
assign reset_logo[26][38] = 9'b100000000;
assign reset_logo[27][1] = 9'b101101101;
assign reset_logo[27][2] = 9'b101101101;
assign reset_logo[27][3] = 9'b101101101;
assign reset_logo[27][4] = 9'b101101101;
assign reset_logo[27][5] = 9'b101101101;
assign reset_logo[27][6] = 9'b101001001;
assign reset_logo[27][7] = 9'b110010001;
assign reset_logo[27][8] = 9'b111101001;
assign reset_logo[27][9] = 9'b111100000;
assign reset_logo[27][10] = 9'b111100100;
assign reset_logo[27][11] = 9'b111100100;
assign reset_logo[27][12] = 9'b111100100;
assign reset_logo[27][13] = 9'b111100100;
assign reset_logo[27][14] = 9'b111100100;
assign reset_logo[27][15] = 9'b111100100;
assign reset_logo[27][16] = 9'b111100100;
assign reset_logo[27][17] = 9'b111100100;
assign reset_logo[27][18] = 9'b111100100;
assign reset_logo[27][19] = 9'b111100100;
assign reset_logo[27][20] = 9'b111100100;
assign reset_logo[27][21] = 9'b111100100;
assign reset_logo[27][22] = 9'b111100100;
assign reset_logo[27][23] = 9'b111100100;
assign reset_logo[27][24] = 9'b111100100;
assign reset_logo[27][25] = 9'b111100100;
assign reset_logo[27][26] = 9'b111100100;
assign reset_logo[27][27] = 9'b111100100;
assign reset_logo[27][28] = 9'b111100100;
assign reset_logo[27][29] = 9'b111100100;
assign reset_logo[27][30] = 9'b111100100;
assign reset_logo[27][31] = 9'b111100100;
assign reset_logo[27][32] = 9'b110001101;
assign reset_logo[27][33] = 9'b101101101;
assign reset_logo[27][34] = 9'b101101101;
assign reset_logo[27][35] = 9'b101001001;
assign reset_logo[27][36] = 9'b101001001;
assign reset_logo[27][37] = 9'b100100100;
assign reset_logo[27][38] = 9'b100100100;
assign reset_logo[28][2] = 9'b101101101;
assign reset_logo[28][3] = 9'b101101101;
assign reset_logo[28][4] = 9'b101101101;
assign reset_logo[28][5] = 9'b101101101;
assign reset_logo[28][6] = 9'b101101001;
assign reset_logo[28][7] = 9'b101001101;
assign reset_logo[28][8] = 9'b110110001;
assign reset_logo[28][9] = 9'b111100100;
assign reset_logo[28][10] = 9'b111100000;
assign reset_logo[28][11] = 9'b111100100;
assign reset_logo[28][12] = 9'b111100100;
assign reset_logo[28][13] = 9'b111100100;
assign reset_logo[28][14] = 9'b111100100;
assign reset_logo[28][15] = 9'b111100100;
assign reset_logo[28][16] = 9'b111100100;
assign reset_logo[28][17] = 9'b111100100;
assign reset_logo[28][18] = 9'b111100100;
assign reset_logo[28][19] = 9'b111100100;
assign reset_logo[28][20] = 9'b111100100;
assign reset_logo[28][21] = 9'b111100100;
assign reset_logo[28][22] = 9'b111100100;
assign reset_logo[28][23] = 9'b111100100;
assign reset_logo[28][24] = 9'b111100100;
assign reset_logo[28][25] = 9'b111100100;
assign reset_logo[28][26] = 9'b111100100;
assign reset_logo[28][27] = 9'b111100100;
assign reset_logo[28][28] = 9'b111100100;
assign reset_logo[28][29] = 9'b111100100;
assign reset_logo[28][30] = 9'b111100100;
assign reset_logo[28][31] = 9'b111101101;
assign reset_logo[28][32] = 9'b101110001;
assign reset_logo[28][33] = 9'b101101101;
assign reset_logo[28][34] = 9'b101101101;
assign reset_logo[28][35] = 9'b101101101;
assign reset_logo[28][36] = 9'b101001000;
assign reset_logo[28][37] = 9'b100100100;
assign reset_logo[29][2] = 9'b101101101;
assign reset_logo[29][3] = 9'b101101101;
assign reset_logo[29][4] = 9'b101101101;
assign reset_logo[29][5] = 9'b101101101;
assign reset_logo[29][6] = 9'b101101001;
assign reset_logo[29][7] = 9'b101001000;
assign reset_logo[29][8] = 9'b101101101;
assign reset_logo[29][9] = 9'b111110001;
assign reset_logo[29][10] = 9'b111100100;
assign reset_logo[29][11] = 9'b111100000;
assign reset_logo[29][12] = 9'b111100100;
assign reset_logo[29][13] = 9'b111100100;
assign reset_logo[29][14] = 9'b111100100;
assign reset_logo[29][15] = 9'b111100100;
assign reset_logo[29][16] = 9'b111100100;
assign reset_logo[29][17] = 9'b111100100;
assign reset_logo[29][18] = 9'b111100100;
assign reset_logo[29][19] = 9'b111100100;
assign reset_logo[29][20] = 9'b111100100;
assign reset_logo[29][21] = 9'b111100100;
assign reset_logo[29][22] = 9'b111100100;
assign reset_logo[29][23] = 9'b111100100;
assign reset_logo[29][24] = 9'b111100100;
assign reset_logo[29][25] = 9'b111100100;
assign reset_logo[29][26] = 9'b111100100;
assign reset_logo[29][27] = 9'b111100100;
assign reset_logo[29][28] = 9'b111100100;
assign reset_logo[29][29] = 9'b111100100;
assign reset_logo[29][30] = 9'b111101101;
assign reset_logo[29][31] = 9'b110010001;
assign reset_logo[29][32] = 9'b110010001;
assign reset_logo[29][33] = 9'b110001101;
assign reset_logo[29][34] = 9'b101101101;
assign reset_logo[29][35] = 9'b101001001;
assign reset_logo[29][36] = 9'b101001000;
assign reset_logo[29][37] = 9'b100100100;
assign reset_logo[30][3] = 9'b101101101;
assign reset_logo[30][4] = 9'b101101101;
assign reset_logo[30][5] = 9'b101101101;
assign reset_logo[30][6] = 9'b101101101;
assign reset_logo[30][7] = 9'b101001001;
assign reset_logo[30][8] = 9'b101001000;
assign reset_logo[30][9] = 9'b101101101;
assign reset_logo[30][10] = 9'b111110001;
assign reset_logo[30][11] = 9'b111100100;
assign reset_logo[30][12] = 9'b111100000;
assign reset_logo[30][13] = 9'b111100000;
assign reset_logo[30][14] = 9'b111100100;
assign reset_logo[30][15] = 9'b111100100;
assign reset_logo[30][16] = 9'b111100100;
assign reset_logo[30][17] = 9'b111100100;
assign reset_logo[30][18] = 9'b111100100;
assign reset_logo[30][19] = 9'b111100100;
assign reset_logo[30][20] = 9'b111100100;
assign reset_logo[30][21] = 9'b111100100;
assign reset_logo[30][22] = 9'b111100100;
assign reset_logo[30][23] = 9'b111100100;
assign reset_logo[30][24] = 9'b111100100;
assign reset_logo[30][25] = 9'b111100100;
assign reset_logo[30][26] = 9'b111100100;
assign reset_logo[30][27] = 9'b111100000;
assign reset_logo[30][28] = 9'b111100100;
assign reset_logo[30][29] = 9'b111101101;
assign reset_logo[30][30] = 9'b110110101;
assign reset_logo[30][31] = 9'b110010001;
assign reset_logo[30][32] = 9'b110010001;
assign reset_logo[30][33] = 9'b110010001;
assign reset_logo[30][34] = 9'b101101101;
assign reset_logo[30][35] = 9'b101001001;
assign reset_logo[30][36] = 9'b100100100;
assign reset_logo[31][4] = 9'b101101101;
assign reset_logo[31][5] = 9'b101001001;
assign reset_logo[31][6] = 9'b101101101;
assign reset_logo[31][7] = 9'b101001001;
assign reset_logo[31][8] = 9'b101001001;
assign reset_logo[31][9] = 9'b101001000;
assign reset_logo[31][10] = 9'b101001101;
assign reset_logo[31][11] = 9'b110010001;
assign reset_logo[31][12] = 9'b111101001;
assign reset_logo[31][13] = 9'b111100000;
assign reset_logo[31][14] = 9'b111100000;
assign reset_logo[31][15] = 9'b111100000;
assign reset_logo[31][16] = 9'b111100100;
assign reset_logo[31][17] = 9'b111100100;
assign reset_logo[31][18] = 9'b111100100;
assign reset_logo[31][19] = 9'b111100100;
assign reset_logo[31][20] = 9'b111100100;
assign reset_logo[31][21] = 9'b111100100;
assign reset_logo[31][22] = 9'b111100100;
assign reset_logo[31][23] = 9'b111100100;
assign reset_logo[31][24] = 9'b111100100;
assign reset_logo[31][25] = 9'b111100000;
assign reset_logo[31][26] = 9'b111100000;
assign reset_logo[31][27] = 9'b111101000;
assign reset_logo[31][28] = 9'b111110001;
assign reset_logo[31][29] = 9'b110010001;
assign reset_logo[31][30] = 9'b110010001;
assign reset_logo[31][31] = 9'b110110010;
assign reset_logo[31][32] = 9'b110010001;
assign reset_logo[31][33] = 9'b110010001;
assign reset_logo[31][34] = 9'b101101101;
assign reset_logo[31][35] = 9'b101001001;
assign reset_logo[31][36] = 9'b100100100;
assign reset_logo[32][4] = 9'b101101101;
assign reset_logo[32][5] = 9'b101101101;
assign reset_logo[32][6] = 9'b101001001;
assign reset_logo[32][7] = 9'b101101101;
assign reset_logo[32][8] = 9'b101001001;
assign reset_logo[32][9] = 9'b101001000;
assign reset_logo[32][10] = 9'b101001000;
assign reset_logo[32][11] = 9'b101001000;
assign reset_logo[32][12] = 9'b101101101;
assign reset_logo[32][13] = 9'b111110001;
assign reset_logo[32][14] = 9'b111101001;
assign reset_logo[32][15] = 9'b111100100;
assign reset_logo[32][16] = 9'b111100000;
assign reset_logo[32][17] = 9'b111100000;
assign reset_logo[32][18] = 9'b111100000;
assign reset_logo[32][19] = 9'b111100000;
assign reset_logo[32][20] = 9'b111100000;
assign reset_logo[32][21] = 9'b111100000;
assign reset_logo[32][22] = 9'b111100000;
assign reset_logo[32][23] = 9'b111100000;
assign reset_logo[32][24] = 9'b111100100;
assign reset_logo[32][25] = 9'b111101000;
assign reset_logo[32][26] = 9'b111101101;
assign reset_logo[32][27] = 9'b110010001;
assign reset_logo[32][28] = 9'b101110001;
assign reset_logo[32][29] = 9'b110010001;
assign reset_logo[32][30] = 9'b110010001;
assign reset_logo[32][31] = 9'b110010001;
assign reset_logo[32][32] = 9'b110010010;
assign reset_logo[32][33] = 9'b101101101;
assign reset_logo[32][34] = 9'b101001001;
assign reset_logo[32][35] = 9'b101001000;
assign reset_logo[33][5] = 9'b101101101;
assign reset_logo[33][6] = 9'b101001001;
assign reset_logo[33][7] = 9'b101001001;
assign reset_logo[33][8] = 9'b101101101;
assign reset_logo[33][9] = 9'b101001001;
assign reset_logo[33][10] = 9'b101001000;
assign reset_logo[33][11] = 9'b101001000;
assign reset_logo[33][12] = 9'b100100100;
assign reset_logo[33][13] = 9'b101001001;
assign reset_logo[33][14] = 9'b101101101;
assign reset_logo[33][15] = 9'b110110001;
assign reset_logo[33][16] = 9'b111101101;
assign reset_logo[33][17] = 9'b111101001;
assign reset_logo[33][18] = 9'b111101000;
assign reset_logo[33][19] = 9'b111100100;
assign reset_logo[33][20] = 9'b111100100;
assign reset_logo[33][21] = 9'b111101000;
assign reset_logo[33][22] = 9'b111101001;
assign reset_logo[33][23] = 9'b111101101;
assign reset_logo[33][24] = 9'b110101101;
assign reset_logo[33][25] = 9'b110001101;
assign reset_logo[33][26] = 9'b101101101;
assign reset_logo[33][27] = 9'b101101101;
assign reset_logo[33][28] = 9'b101101101;
assign reset_logo[33][29] = 9'b110001101;
assign reset_logo[33][30] = 9'b110010001;
assign reset_logo[33][31] = 9'b110010001;
assign reset_logo[33][32] = 9'b101101101;
assign reset_logo[33][33] = 9'b101101101;
assign reset_logo[33][34] = 9'b101001001;
assign reset_logo[34][6] = 9'b101001001;
assign reset_logo[34][7] = 9'b101001001;
assign reset_logo[34][8] = 9'b101001001;
assign reset_logo[34][9] = 9'b101001001;
assign reset_logo[34][10] = 9'b101001001;
assign reset_logo[34][11] = 9'b101001000;
assign reset_logo[34][12] = 9'b100100100;
assign reset_logo[34][13] = 9'b100100100;
assign reset_logo[34][14] = 9'b100100100;
assign reset_logo[34][15] = 9'b100100100;
assign reset_logo[34][16] = 9'b101001001;
assign reset_logo[34][17] = 9'b101101101;
assign reset_logo[34][18] = 9'b101101101;
assign reset_logo[34][19] = 9'b101101101;
assign reset_logo[34][20] = 9'b110001101;
assign reset_logo[34][21] = 9'b101101101;
assign reset_logo[34][22] = 9'b101101101;
assign reset_logo[34][23] = 9'b101001101;
assign reset_logo[34][24] = 9'b101001001;
assign reset_logo[34][25] = 9'b101001001;
assign reset_logo[34][26] = 9'b101101101;
assign reset_logo[34][27] = 9'b101101101;
assign reset_logo[34][28] = 9'b101101101;
assign reset_logo[34][29] = 9'b101101101;
assign reset_logo[34][30] = 9'b101101101;
assign reset_logo[34][31] = 9'b101101101;
assign reset_logo[34][32] = 9'b101001001;
assign reset_logo[34][33] = 9'b101001001;
assign reset_logo[35][7] = 9'b101001001;
assign reset_logo[35][8] = 9'b101001001;
assign reset_logo[35][9] = 9'b101001000;
assign reset_logo[35][10] = 9'b101001001;
assign reset_logo[35][11] = 9'b101001001;
assign reset_logo[35][12] = 9'b100100100;
assign reset_logo[35][13] = 9'b100100100;
assign reset_logo[35][14] = 9'b100100100;
assign reset_logo[35][15] = 9'b100100000;
assign reset_logo[35][16] = 9'b100100100;
assign reset_logo[35][17] = 9'b100100100;
assign reset_logo[35][18] = 9'b100100100;
assign reset_logo[35][19] = 9'b100100100;
assign reset_logo[35][20] = 9'b100100100;
assign reset_logo[35][21] = 9'b100100100;
assign reset_logo[35][22] = 9'b101001000;
assign reset_logo[35][23] = 9'b101001000;
assign reset_logo[35][24] = 9'b101001000;
assign reset_logo[35][25] = 9'b101001001;
assign reset_logo[35][26] = 9'b101001001;
assign reset_logo[35][27] = 9'b101001001;
assign reset_logo[35][28] = 9'b101101101;
assign reset_logo[35][29] = 9'b101001001;
assign reset_logo[35][30] = 9'b101001001;
assign reset_logo[35][31] = 9'b101001001;
assign reset_logo[35][32] = 9'b101001000;
assign reset_logo[36][8] = 9'b101001000;
assign reset_logo[36][9] = 9'b101001000;
assign reset_logo[36][10] = 9'b101001000;
assign reset_logo[36][11] = 9'b100100100;
assign reset_logo[36][12] = 9'b100100100;
assign reset_logo[36][13] = 9'b100100100;
assign reset_logo[36][14] = 9'b100100100;
assign reset_logo[36][15] = 9'b100000100;
assign reset_logo[36][16] = 9'b100000000;
assign reset_logo[36][17] = 9'b100000000;
assign reset_logo[36][18] = 9'b100100000;
assign reset_logo[36][19] = 9'b100100100;
assign reset_logo[36][20] = 9'b100100100;
assign reset_logo[36][21] = 9'b100100100;
assign reset_logo[36][22] = 9'b100100100;
assign reset_logo[36][23] = 9'b100100100;
assign reset_logo[36][24] = 9'b100100100;
assign reset_logo[36][25] = 9'b101001000;
assign reset_logo[36][26] = 9'b101001001;
assign reset_logo[36][27] = 9'b101001001;
assign reset_logo[36][28] = 9'b101001000;
assign reset_logo[36][29] = 9'b101001000;
assign reset_logo[36][30] = 9'b100100100;
assign reset_logo[36][31] = 9'b100100100;
assign reset_logo[37][10] = 9'b101001000;
assign reset_logo[37][11] = 9'b100100100;
assign reset_logo[37][12] = 9'b100100100;
assign reset_logo[37][13] = 9'b100100100;
assign reset_logo[37][14] = 9'b100100100;
assign reset_logo[37][15] = 9'b100100100;
assign reset_logo[37][16] = 9'b100000000;
assign reset_logo[37][17] = 9'b100000000;
assign reset_logo[37][18] = 9'b100000000;
assign reset_logo[37][19] = 9'b100000000;
assign reset_logo[37][20] = 9'b100000000;
assign reset_logo[37][21] = 9'b100100100;
assign reset_logo[37][22] = 9'b100100100;
assign reset_logo[37][23] = 9'b100100100;
assign reset_logo[37][24] = 9'b100100100;
assign reset_logo[37][25] = 9'b100100100;
assign reset_logo[37][26] = 9'b100100100;
assign reset_logo[37][27] = 9'b100100100;
assign reset_logo[37][28] = 9'b100100100;
assign reset_logo[37][29] = 9'b100100100;
assign reset_logo[38][12] = 9'b100100100;
assign reset_logo[38][13] = 9'b100100100;
assign reset_logo[38][14] = 9'b100100100;
assign reset_logo[38][15] = 9'b100100100;
assign reset_logo[38][16] = 9'b100000000;
assign reset_logo[38][17] = 9'b100000000;
assign reset_logo[38][18] = 9'b100000000;
assign reset_logo[38][19] = 9'b100000000;
assign reset_logo[38][20] = 9'b100000000;
assign reset_logo[38][21] = 9'b100000000;
assign reset_logo[38][22] = 9'b100000000;
assign reset_logo[38][23] = 9'b100000000;
assign reset_logo[38][24] = 9'b100000000;
assign reset_logo[38][25] = 9'b100000000;
assign reset_logo[38][26] = 9'b100100100;
assign reset_logo[38][27] = 9'b100100100;
assign reset_logo[39][15] = 9'b100000000;
assign reset_logo[39][16] = 9'b100000000;
assign reset_logo[39][17] = 9'b100000000;
assign reset_logo[39][18] = 9'b100000000;
assign reset_logo[39][19] = 9'b100000000;
assign reset_logo[39][20] = 9'b100000000;
assign reset_logo[39][21] = 9'b100000000;
assign reset_logo[39][22] = 9'b100000000;
assign reset_logo[39][23] = 9'b100000000;
assign reset_logo[39][24] = 9'b100000000;
//Total de Lineas = 1279
endmodule

