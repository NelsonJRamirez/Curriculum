`timescale 1ns / 1ps
module logo_start (
input enable,
input clock,
input [9:0] posx, posy,
input [9:0] hcount,
input [9:0] vcount,
output reg[2:0] red,
output reg[2:0] green,
output reg[1:0] blue,
output reg data);

always @(posedge clock)
begin
	if(enable)
	begin
		if(hcount >= posx & hcount < posx + RESOLUCION_X & vcount >= posy & vcount < posy + RESOLUCION_Y)
		begin
			if (logo_start[vcount - posy][hcount - posx][8] == 1'b1)
			begin
				red   <= logo_start[vcount- posy][hcount- posx][7:5];
				green <= logo_start[vcount- posy][hcount- posx][4:2];
            blue 	<= logo_start[vcount- posy][hcount- posx][1:0];
				data  <= 1'b1;
			end
			else
				data <= 0;
			end
		else
		data <= 0;
	end
end

parameter RESOLUCION_X = 40;
parameter RESOLUCION_Y = 20;
wire [8:0] logo_start[RESOLUCION_Y - 1'b1 : 0][RESOLUCION_X - 1'b1 : 0];
assign logo_start[1][5] = 9'b100000000;
assign logo_start[1][6] = 9'b100000000;
assign logo_start[1][7] = 9'b100000000;
assign logo_start[1][8] = 9'b100000000;
assign logo_start[1][9] = 9'b100000000;
assign logo_start[1][10] = 9'b100000000;
assign logo_start[1][11] = 9'b100000000;
assign logo_start[1][12] = 9'b100000000;
assign logo_start[1][13] = 9'b100000000;
assign logo_start[1][14] = 9'b100000000;
assign logo_start[1][15] = 9'b100000000;
assign logo_start[1][16] = 9'b100000000;
assign logo_start[1][17] = 9'b100000000;
assign logo_start[1][18] = 9'b100000000;
assign logo_start[1][19] = 9'b100000000;
assign logo_start[1][20] = 9'b100000000;
assign logo_start[1][21] = 9'b100000000;
assign logo_start[1][22] = 9'b100000000;
assign logo_start[1][23] = 9'b100000000;
assign logo_start[1][24] = 9'b100000000;
assign logo_start[1][25] = 9'b100000000;
assign logo_start[1][26] = 9'b100000000;
assign logo_start[1][27] = 9'b100000000;
assign logo_start[1][28] = 9'b100000000;
assign logo_start[1][29] = 9'b100000000;
assign logo_start[1][30] = 9'b100000000;
assign logo_start[1][31] = 9'b100000000;
assign logo_start[1][32] = 9'b100000000;
assign logo_start[1][33] = 9'b100000000;
assign logo_start[1][34] = 9'b100000000;
assign logo_start[1][35] = 9'b100000000;
assign logo_start[2][3] = 9'b100000000;
assign logo_start[2][4] = 9'b100000000;
assign logo_start[2][5] = 9'b100100000;
assign logo_start[2][6] = 9'b100100000;
assign logo_start[2][7] = 9'b100100000;
assign logo_start[2][8] = 9'b100100000;
assign logo_start[2][9] = 9'b100100000;
assign logo_start[2][10] = 9'b100100000;
assign logo_start[2][11] = 9'b100100000;
assign logo_start[2][12] = 9'b100100000;
assign logo_start[2][13] = 9'b100100000;
assign logo_start[2][14] = 9'b100100000;
assign logo_start[2][15] = 9'b100100000;
assign logo_start[2][16] = 9'b100100000;
assign logo_start[2][17] = 9'b100100000;
assign logo_start[2][18] = 9'b100100000;
assign logo_start[2][19] = 9'b100100000;
assign logo_start[2][20] = 9'b100100000;
assign logo_start[2][21] = 9'b100100000;
assign logo_start[2][22] = 9'b100100000;
assign logo_start[2][23] = 9'b100100000;
assign logo_start[2][24] = 9'b100100000;
assign logo_start[2][25] = 9'b100100000;
assign logo_start[2][26] = 9'b100100000;
assign logo_start[2][27] = 9'b100100000;
assign logo_start[2][28] = 9'b100100000;
assign logo_start[2][29] = 9'b100100000;
assign logo_start[2][30] = 9'b100100000;
assign logo_start[2][31] = 9'b100100000;
assign logo_start[2][32] = 9'b100100000;
assign logo_start[2][33] = 9'b100100000;
assign logo_start[2][34] = 9'b100100000;
assign logo_start[2][35] = 9'b100100000;
assign logo_start[2][36] = 9'b100000000;
assign logo_start[3][2] = 9'b100000000;
assign logo_start[3][3] = 9'b100000000;
assign logo_start[3][4] = 9'b110000000;
assign logo_start[3][5] = 9'b111100100;
assign logo_start[3][6] = 9'b111100100;
assign logo_start[3][7] = 9'b111100100;
assign logo_start[3][8] = 9'b111100100;
assign logo_start[3][9] = 9'b111100100;
assign logo_start[3][10] = 9'b111100100;
assign logo_start[3][11] = 9'b111100100;
assign logo_start[3][12] = 9'b111100100;
assign logo_start[3][13] = 9'b111100100;
assign logo_start[3][14] = 9'b111100100;
assign logo_start[3][15] = 9'b111100100;
assign logo_start[3][16] = 9'b111100100;
assign logo_start[3][17] = 9'b111100100;
assign logo_start[3][18] = 9'b111100100;
assign logo_start[3][19] = 9'b111100100;
assign logo_start[3][20] = 9'b111100100;
assign logo_start[3][21] = 9'b111100100;
assign logo_start[3][22] = 9'b111100000;
assign logo_start[3][23] = 9'b111100000;
assign logo_start[3][24] = 9'b111100000;
assign logo_start[3][25] = 9'b111100000;
assign logo_start[3][26] = 9'b111100000;
assign logo_start[3][27] = 9'b111100000;
assign logo_start[3][28] = 9'b111100000;
assign logo_start[3][29] = 9'b111100000;
assign logo_start[3][30] = 9'b111100000;
assign logo_start[3][31] = 9'b111100000;
assign logo_start[3][32] = 9'b111100000;
assign logo_start[3][33] = 9'b111100000;
assign logo_start[3][34] = 9'b111100000;
assign logo_start[3][35] = 9'b111100000;
assign logo_start[3][36] = 9'b100100000;
assign logo_start[3][37] = 9'b100000000;
assign logo_start[4][2] = 9'b100000000;
assign logo_start[4][3] = 9'b110000000;
assign logo_start[4][4] = 9'b111100100;
assign logo_start[4][5] = 9'b111100100;
assign logo_start[4][6] = 9'b111100100;
assign logo_start[4][7] = 9'b111100100;
assign logo_start[4][8] = 9'b111100100;
assign logo_start[4][9] = 9'b111100100;
assign logo_start[4][10] = 9'b111100100;
assign logo_start[4][11] = 9'b111100100;
assign logo_start[4][12] = 9'b111100100;
assign logo_start[4][13] = 9'b111100100;
assign logo_start[4][14] = 9'b111100100;
assign logo_start[4][15] = 9'b111100100;
assign logo_start[4][16] = 9'b111100100;
assign logo_start[4][17] = 9'b111100100;
assign logo_start[4][18] = 9'b111100100;
assign logo_start[4][19] = 9'b111100100;
assign logo_start[4][20] = 9'b111100000;
assign logo_start[4][21] = 9'b110100000;
assign logo_start[4][22] = 9'b111100000;
assign logo_start[4][23] = 9'b111100000;
assign logo_start[4][24] = 9'b110100000;
assign logo_start[4][25] = 9'b110100000;
assign logo_start[4][26] = 9'b110100000;
assign logo_start[4][27] = 9'b110100000;
assign logo_start[4][28] = 9'b111100000;
assign logo_start[4][29] = 9'b111100000;
assign logo_start[4][30] = 9'b110100000;
assign logo_start[4][31] = 9'b110100000;
assign logo_start[4][32] = 9'b110100000;
assign logo_start[4][33] = 9'b110100000;
assign logo_start[4][34] = 9'b110100000;
assign logo_start[4][35] = 9'b110100000;
assign logo_start[4][36] = 9'b110000000;
assign logo_start[4][37] = 9'b100100000;
assign logo_start[4][38] = 9'b100000000;
assign logo_start[5][2] = 9'b100000000;
assign logo_start[5][3] = 9'b111100100;
assign logo_start[5][4] = 9'b111100100;
assign logo_start[5][5] = 9'b111100000;
assign logo_start[5][6] = 9'b100100000;
assign logo_start[5][7] = 9'b100000000;
assign logo_start[5][8] = 9'b100000000;
assign logo_start[5][9] = 9'b100000000;
assign logo_start[5][10] = 9'b110100000;
assign logo_start[5][11] = 9'b101100000;
assign logo_start[5][12] = 9'b100000000;
assign logo_start[5][13] = 9'b100000000;
assign logo_start[5][14] = 9'b100000000;
assign logo_start[5][15] = 9'b100000000;
assign logo_start[5][16] = 9'b101000000;
assign logo_start[5][17] = 9'b111100100;
assign logo_start[5][18] = 9'b101100000;
assign logo_start[5][19] = 9'b100000000;
assign logo_start[5][20] = 9'b100000000;
assign logo_start[5][21] = 9'b100000000;
assign logo_start[5][22] = 9'b110100000;
assign logo_start[5][23] = 9'b110100000;
assign logo_start[5][24] = 9'b100000000;
assign logo_start[5][25] = 9'b100000000;
assign logo_start[5][26] = 9'b100000000;
assign logo_start[5][27] = 9'b100000000;
assign logo_start[5][28] = 9'b110000000;
assign logo_start[5][29] = 9'b111100000;
assign logo_start[5][30] = 9'b100100000;
assign logo_start[5][31] = 9'b100000000;
assign logo_start[5][32] = 9'b100000000;
assign logo_start[5][33] = 9'b100000000;
assign logo_start[5][34] = 9'b100000000;
assign logo_start[5][35] = 9'b101100000;
assign logo_start[5][36] = 9'b111100000;
assign logo_start[5][37] = 9'b101000000;
assign logo_start[5][38] = 9'b100000000;
assign logo_start[6][2] = 9'b100000000;
assign logo_start[6][3] = 9'b111100000;
assign logo_start[6][4] = 9'b111100100;
assign logo_start[6][5] = 9'b100100000;
assign logo_start[6][6] = 9'b101000000;
assign logo_start[6][7] = 9'b111100000;
assign logo_start[6][8] = 9'b111100000;
assign logo_start[6][9] = 9'b111100000;
assign logo_start[6][10] = 9'b111100100;
assign logo_start[6][11] = 9'b111100100;
assign logo_start[6][12] = 9'b111100000;
assign logo_start[6][13] = 9'b100000000;
assign logo_start[6][14] = 9'b100000000;
assign logo_start[6][15] = 9'b110100000;
assign logo_start[6][16] = 9'b111100100;
assign logo_start[6][17] = 9'b110000000;
assign logo_start[6][18] = 9'b100000000;
assign logo_start[6][19] = 9'b110000000;
assign logo_start[6][20] = 9'b110100000;
assign logo_start[6][21] = 9'b101000000;
assign logo_start[6][22] = 9'b100100000;
assign logo_start[6][23] = 9'b110000000;
assign logo_start[6][24] = 9'b100000000;
assign logo_start[6][25] = 9'b101100000;
assign logo_start[6][26] = 9'b110100000;
assign logo_start[6][27] = 9'b101100000;
assign logo_start[6][28] = 9'b100000000;
assign logo_start[6][29] = 9'b110100000;
assign logo_start[6][30] = 9'b110100000;
assign logo_start[6][31] = 9'b101100000;
assign logo_start[6][32] = 9'b100000000;
assign logo_start[6][33] = 9'b100100000;
assign logo_start[6][34] = 9'b110000000;
assign logo_start[6][35] = 9'b110000000;
assign logo_start[6][36] = 9'b110100000;
assign logo_start[6][37] = 9'b100100000;
assign logo_start[6][38] = 9'b100000000;
assign logo_start[7][2] = 9'b100000000;
assign logo_start[7][3] = 9'b111100000;
assign logo_start[7][4] = 9'b111100100;
assign logo_start[7][5] = 9'b100100000;
assign logo_start[7][6] = 9'b110100000;
assign logo_start[7][7] = 9'b111100100;
assign logo_start[7][8] = 9'b111100100;
assign logo_start[7][9] = 9'b111100100;
assign logo_start[7][10] = 9'b111100100;
assign logo_start[7][11] = 9'b111100100;
assign logo_start[7][12] = 9'b111100100;
assign logo_start[7][13] = 9'b101100000;
assign logo_start[7][14] = 9'b101000000;
assign logo_start[7][15] = 9'b111100100;
assign logo_start[7][16] = 9'b111100100;
assign logo_start[7][17] = 9'b110000000;
assign logo_start[7][18] = 9'b100100000;
assign logo_start[7][19] = 9'b111100100;
assign logo_start[7][20] = 9'b111100000;
assign logo_start[7][21] = 9'b110000000;
assign logo_start[7][22] = 9'b100000000;
assign logo_start[7][23] = 9'b110000000;
assign logo_start[7][24] = 9'b100000000;
assign logo_start[7][25] = 9'b111100000;
assign logo_start[7][26] = 9'b111100000;
assign logo_start[7][27] = 9'b111100000;
assign logo_start[7][28] = 9'b100000000;
assign logo_start[7][29] = 9'b110000000;
assign logo_start[7][30] = 9'b111100000;
assign logo_start[7][31] = 9'b111100000;
assign logo_start[7][32] = 9'b100100000;
assign logo_start[7][33] = 9'b101100000;
assign logo_start[7][34] = 9'b110100000;
assign logo_start[7][35] = 9'b110000000;
assign logo_start[7][36] = 9'b110100000;
assign logo_start[7][37] = 9'b100100000;
assign logo_start[7][38] = 9'b100000000;
assign logo_start[8][2] = 9'b100000000;
assign logo_start[8][3] = 9'b111100000;
assign logo_start[8][4] = 9'b111100100;
assign logo_start[8][5] = 9'b100000000;
assign logo_start[8][6] = 9'b110000000;
assign logo_start[8][7] = 9'b111100100;
assign logo_start[8][8] = 9'b111100100;
assign logo_start[8][9] = 9'b111100100;
assign logo_start[8][10] = 9'b111100100;
assign logo_start[8][11] = 9'b111100100;
assign logo_start[8][12] = 9'b111100100;
assign logo_start[8][13] = 9'b101000000;
assign logo_start[8][14] = 9'b101000000;
assign logo_start[8][15] = 9'b111100100;
assign logo_start[8][16] = 9'b111100100;
assign logo_start[8][17] = 9'b101100000;
assign logo_start[8][18] = 9'b100100000;
assign logo_start[8][19] = 9'b111100000;
assign logo_start[8][20] = 9'b111100100;
assign logo_start[8][21] = 9'b110000000;
assign logo_start[8][22] = 9'b100000000;
assign logo_start[8][23] = 9'b110000000;
assign logo_start[8][24] = 9'b100000000;
assign logo_start[8][25] = 9'b110100000;
assign logo_start[8][26] = 9'b111100100;
assign logo_start[8][27] = 9'b110100000;
assign logo_start[8][28] = 9'b100000000;
assign logo_start[8][29] = 9'b110000000;
assign logo_start[8][30] = 9'b111100000;
assign logo_start[8][31] = 9'b110100000;
assign logo_start[8][32] = 9'b100000000;
assign logo_start[8][33] = 9'b101100000;
assign logo_start[8][34] = 9'b110100000;
assign logo_start[8][35] = 9'b110000000;
assign logo_start[8][36] = 9'b110100000;
assign logo_start[8][37] = 9'b100100000;
assign logo_start[8][38] = 9'b100000000;
assign logo_start[9][2] = 9'b100000000;
assign logo_start[9][3] = 9'b111100000;
assign logo_start[9][4] = 9'b111100100;
assign logo_start[9][5] = 9'b101100000;
assign logo_start[9][6] = 9'b100000000;
assign logo_start[9][7] = 9'b101000000;
assign logo_start[9][8] = 9'b101000000;
assign logo_start[9][9] = 9'b110100000;
assign logo_start[9][10] = 9'b111100100;
assign logo_start[9][11] = 9'b111100100;
assign logo_start[9][12] = 9'b111100100;
assign logo_start[9][13] = 9'b101000000;
assign logo_start[9][14] = 9'b101000000;
assign logo_start[9][15] = 9'b111100100;
assign logo_start[9][16] = 9'b111100100;
assign logo_start[9][17] = 9'b101100000;
assign logo_start[9][18] = 9'b100000000;
assign logo_start[9][19] = 9'b100100000;
assign logo_start[9][20] = 9'b101000000;
assign logo_start[9][21] = 9'b100000000;
assign logo_start[9][22] = 9'b100100000;
assign logo_start[9][23] = 9'b110000000;
assign logo_start[9][24] = 9'b100000000;
assign logo_start[9][25] = 9'b100100000;
assign logo_start[9][26] = 9'b101000000;
assign logo_start[9][27] = 9'b100100000;
assign logo_start[9][28] = 9'b101100000;
assign logo_start[9][29] = 9'b111100000;
assign logo_start[9][30] = 9'b110100000;
assign logo_start[9][31] = 9'b110000000;
assign logo_start[9][32] = 9'b100000000;
assign logo_start[9][33] = 9'b101100000;
assign logo_start[9][34] = 9'b110100000;
assign logo_start[9][35] = 9'b110000000;
assign logo_start[9][36] = 9'b110100000;
assign logo_start[9][37] = 9'b100100000;
assign logo_start[9][38] = 9'b100000000;
assign logo_start[10][2] = 9'b100000000;
assign logo_start[10][3] = 9'b111100000;
assign logo_start[10][4] = 9'b111100100;
assign logo_start[10][5] = 9'b111100100;
assign logo_start[10][6] = 9'b101100000;
assign logo_start[10][7] = 9'b101000000;
assign logo_start[10][8] = 9'b100100000;
assign logo_start[10][9] = 9'b100000000;
assign logo_start[10][10] = 9'b111100000;
assign logo_start[10][11] = 9'b111100100;
assign logo_start[10][12] = 9'b111100100;
assign logo_start[10][13] = 9'b101000000;
assign logo_start[10][14] = 9'b101000000;
assign logo_start[10][15] = 9'b111100100;
assign logo_start[10][16] = 9'b111100000;
assign logo_start[10][17] = 9'b101100000;
assign logo_start[10][18] = 9'b100000000;
assign logo_start[10][19] = 9'b100100000;
assign logo_start[10][20] = 9'b101000000;
assign logo_start[10][21] = 9'b100000000;
assign logo_start[10][22] = 9'b100100000;
assign logo_start[10][23] = 9'b110000000;
assign logo_start[10][24] = 9'b100000000;
assign logo_start[10][25] = 9'b100100000;
assign logo_start[10][26] = 9'b101000000;
assign logo_start[10][27] = 9'b100100000;
assign logo_start[10][28] = 9'b101100000;
assign logo_start[10][29] = 9'b110100000;
assign logo_start[10][30] = 9'b110000000;
assign logo_start[10][31] = 9'b110000000;
assign logo_start[10][32] = 9'b100000000;
assign logo_start[10][33] = 9'b101100000;
assign logo_start[10][34] = 9'b110100000;
assign logo_start[10][35] = 9'b110000000;
assign logo_start[10][36] = 9'b110100000;
assign logo_start[10][37] = 9'b100100000;
assign logo_start[10][38] = 9'b100000000;
assign logo_start[11][2] = 9'b100000000;
assign logo_start[11][3] = 9'b111100000;
assign logo_start[11][4] = 9'b111100100;
assign logo_start[11][5] = 9'b111100100;
assign logo_start[11][6] = 9'b111100100;
assign logo_start[11][7] = 9'b111100100;
assign logo_start[11][8] = 9'b111100100;
assign logo_start[11][9] = 9'b100100000;
assign logo_start[11][10] = 9'b101100000;
assign logo_start[11][11] = 9'b111100100;
assign logo_start[11][12] = 9'b111100100;
assign logo_start[11][13] = 9'b101100000;
assign logo_start[11][14] = 9'b100100000;
assign logo_start[11][15] = 9'b111100000;
assign logo_start[11][16] = 9'b111100000;
assign logo_start[11][17] = 9'b101100000;
assign logo_start[11][18] = 9'b100100000;
assign logo_start[11][19] = 9'b111100000;
assign logo_start[11][20] = 9'b111100100;
assign logo_start[11][21] = 9'b110000000;
assign logo_start[11][22] = 9'b100000000;
assign logo_start[11][23] = 9'b110000000;
assign logo_start[11][24] = 9'b100000000;
assign logo_start[11][25] = 9'b110100000;
assign logo_start[11][26] = 9'b111100100;
assign logo_start[11][27] = 9'b110100000;
assign logo_start[11][28] = 9'b100000000;
assign logo_start[11][29] = 9'b101100000;
assign logo_start[11][30] = 9'b110100000;
assign logo_start[11][31] = 9'b110000000;
assign logo_start[11][32] = 9'b100000000;
assign logo_start[11][33] = 9'b101100000;
assign logo_start[11][34] = 9'b110100000;
assign logo_start[11][35] = 9'b110000000;
assign logo_start[11][36] = 9'b110100000;
assign logo_start[11][37] = 9'b100100000;
assign logo_start[11][38] = 9'b100000000;
assign logo_start[12][2] = 9'b100000000;
assign logo_start[12][3] = 9'b111100000;
assign logo_start[12][4] = 9'b111100100;
assign logo_start[12][5] = 9'b111100100;
assign logo_start[12][6] = 9'b111100100;
assign logo_start[12][7] = 9'b111100100;
assign logo_start[12][8] = 9'b111100100;
assign logo_start[12][9] = 9'b101000000;
assign logo_start[12][10] = 9'b101100000;
assign logo_start[12][11] = 9'b111100100;
assign logo_start[12][12] = 9'b111100100;
assign logo_start[12][13] = 9'b101000000;
assign logo_start[12][14] = 9'b101000000;
assign logo_start[12][15] = 9'b111100000;
assign logo_start[12][16] = 9'b111100000;
assign logo_start[12][17] = 9'b101100000;
assign logo_start[12][18] = 9'b100100000;
assign logo_start[12][19] = 9'b111100000;
assign logo_start[12][20] = 9'b111100000;
assign logo_start[12][21] = 9'b110000000;
assign logo_start[12][22] = 9'b100100000;
assign logo_start[12][23] = 9'b110000000;
assign logo_start[12][24] = 9'b100000000;
assign logo_start[12][25] = 9'b111100000;
assign logo_start[12][26] = 9'b111100000;
assign logo_start[12][27] = 9'b110100000;
assign logo_start[12][28] = 9'b100000000;
assign logo_start[12][29] = 9'b110000000;
assign logo_start[12][30] = 9'b110100000;
assign logo_start[12][31] = 9'b110000000;
assign logo_start[12][32] = 9'b100000000;
assign logo_start[12][33] = 9'b101100000;
assign logo_start[12][34] = 9'b110100000;
assign logo_start[12][35] = 9'b110000000;
assign logo_start[12][36] = 9'b110100000;
assign logo_start[12][37] = 9'b100100000;
assign logo_start[12][38] = 9'b100000000;
assign logo_start[13][2] = 9'b100000000;
assign logo_start[13][3] = 9'b111100000;
assign logo_start[13][4] = 9'b111100100;
assign logo_start[13][5] = 9'b111100000;
assign logo_start[13][6] = 9'b111100000;
assign logo_start[13][7] = 9'b111100000;
assign logo_start[13][8] = 9'b110100000;
assign logo_start[13][9] = 9'b100000000;
assign logo_start[13][10] = 9'b110000000;
assign logo_start[13][11] = 9'b111100100;
assign logo_start[13][12] = 9'b111100100;
assign logo_start[13][13] = 9'b101000000;
assign logo_start[13][14] = 9'b101000000;
assign logo_start[13][15] = 9'b111100000;
assign logo_start[13][16] = 9'b111100000;
assign logo_start[13][17] = 9'b101100000;
assign logo_start[13][18] = 9'b100100000;
assign logo_start[13][19] = 9'b111100000;
assign logo_start[13][20] = 9'b111100000;
assign logo_start[13][21] = 9'b110000000;
assign logo_start[13][22] = 9'b100000000;
assign logo_start[13][23] = 9'b110000000;
assign logo_start[13][24] = 9'b100000000;
assign logo_start[13][25] = 9'b111100000;
assign logo_start[13][26] = 9'b111100000;
assign logo_start[13][27] = 9'b110000000;
assign logo_start[13][28] = 9'b100000000;
assign logo_start[13][29] = 9'b110000000;
assign logo_start[13][30] = 9'b110100000;
assign logo_start[13][31] = 9'b110000000;
assign logo_start[13][32] = 9'b100000000;
assign logo_start[13][33] = 9'b101100000;
assign logo_start[13][34] = 9'b110100000;
assign logo_start[13][35] = 9'b110000000;
assign logo_start[13][36] = 9'b110100000;
assign logo_start[13][37] = 9'b100100000;
assign logo_start[13][38] = 9'b100000000;
assign logo_start[14][2] = 9'b100000000;
assign logo_start[14][3] = 9'b111100100;
assign logo_start[14][4] = 9'b111100100;
assign logo_start[14][5] = 9'b100100000;
assign logo_start[14][6] = 9'b100000000;
assign logo_start[14][7] = 9'b100000000;
assign logo_start[14][8] = 9'b100000000;
assign logo_start[14][9] = 9'b101100000;
assign logo_start[14][10] = 9'b111100100;
assign logo_start[14][11] = 9'b111100000;
assign logo_start[14][12] = 9'b111100000;
assign logo_start[14][13] = 9'b101000000;
assign logo_start[14][14] = 9'b101000000;
assign logo_start[14][15] = 9'b111100000;
assign logo_start[14][16] = 9'b111100000;
assign logo_start[14][17] = 9'b101100000;
assign logo_start[14][18] = 9'b100100000;
assign logo_start[14][19] = 9'b111100000;
assign logo_start[14][20] = 9'b111100000;
assign logo_start[14][21] = 9'b110000000;
assign logo_start[14][22] = 9'b100100000;
assign logo_start[14][23] = 9'b110000000;
assign logo_start[14][24] = 9'b100100000;
assign logo_start[14][25] = 9'b110100000;
assign logo_start[14][26] = 9'b110100000;
assign logo_start[14][27] = 9'b110000000;
assign logo_start[14][28] = 9'b100000000;
assign logo_start[14][29] = 9'b110000000;
assign logo_start[14][30] = 9'b110100000;
assign logo_start[14][31] = 9'b110000000;
assign logo_start[14][32] = 9'b100100000;
assign logo_start[14][33] = 9'b101100000;
assign logo_start[14][34] = 9'b110100000;
assign logo_start[14][35] = 9'b110000000;
assign logo_start[14][36] = 9'b110100000;
assign logo_start[14][37] = 9'b101000000;
assign logo_start[14][38] = 9'b100000000;
assign logo_start[15][2] = 9'b100000000;
assign logo_start[15][3] = 9'b110000000;
assign logo_start[15][4] = 9'b111100100;
assign logo_start[15][5] = 9'b111100100;
assign logo_start[15][6] = 9'b111100100;
assign logo_start[15][7] = 9'b111100100;
assign logo_start[15][8] = 9'b111100100;
assign logo_start[15][9] = 9'b111100100;
assign logo_start[15][10] = 9'b111100100;
assign logo_start[15][11] = 9'b111100000;
assign logo_start[15][12] = 9'b111100000;
assign logo_start[15][13] = 9'b111100000;
assign logo_start[15][14] = 9'b111100000;
assign logo_start[15][15] = 9'b111100000;
assign logo_start[15][16] = 9'b111100000;
assign logo_start[15][17] = 9'b111100000;
assign logo_start[15][18] = 9'b110100000;
assign logo_start[15][19] = 9'b111100000;
assign logo_start[15][20] = 9'b111100000;
assign logo_start[15][21] = 9'b111100000;
assign logo_start[15][22] = 9'b110100000;
assign logo_start[15][23] = 9'b111100000;
assign logo_start[15][24] = 9'b110100000;
assign logo_start[15][25] = 9'b110000000;
assign logo_start[15][26] = 9'b110000000;
assign logo_start[15][27] = 9'b110000000;
assign logo_start[15][28] = 9'b110000000;
assign logo_start[15][29] = 9'b110000000;
assign logo_start[15][30] = 9'b110000000;
assign logo_start[15][31] = 9'b110000000;
assign logo_start[15][32] = 9'b110000000;
assign logo_start[15][33] = 9'b110000000;
assign logo_start[15][34] = 9'b110000000;
assign logo_start[15][35] = 9'b110100000;
assign logo_start[15][36] = 9'b110000000;
assign logo_start[15][37] = 9'b100100000;
assign logo_start[15][38] = 9'b100000000;
assign logo_start[16][2] = 9'b100000000;
assign logo_start[16][3] = 9'b100000000;
assign logo_start[16][4] = 9'b110000000;
assign logo_start[16][5] = 9'b111100100;
assign logo_start[16][6] = 9'b111100100;
assign logo_start[16][7] = 9'b111100100;
assign logo_start[16][8] = 9'b111100100;
assign logo_start[16][9] = 9'b111100100;
assign logo_start[16][10] = 9'b111100000;
assign logo_start[16][11] = 9'b111100000;
assign logo_start[16][12] = 9'b111100000;
assign logo_start[16][13] = 9'b111100000;
assign logo_start[16][14] = 9'b111100000;
assign logo_start[16][15] = 9'b111100000;
assign logo_start[16][16] = 9'b111100000;
assign logo_start[16][17] = 9'b111100000;
assign logo_start[16][18] = 9'b111100000;
assign logo_start[16][19] = 9'b111100000;
assign logo_start[16][20] = 9'b111100000;
assign logo_start[16][21] = 9'b111100000;
assign logo_start[16][22] = 9'b111100000;
assign logo_start[16][23] = 9'b111100000;
assign logo_start[16][24] = 9'b110100000;
assign logo_start[16][25] = 9'b110000000;
assign logo_start[16][26] = 9'b110000000;
assign logo_start[16][27] = 9'b110100000;
assign logo_start[16][28] = 9'b110100000;
assign logo_start[16][29] = 9'b110100000;
assign logo_start[16][30] = 9'b110100000;
assign logo_start[16][31] = 9'b110100000;
assign logo_start[16][32] = 9'b110100000;
assign logo_start[16][33] = 9'b110100000;
assign logo_start[16][34] = 9'b110100000;
assign logo_start[16][35] = 9'b110000000;
assign logo_start[16][36] = 9'b100100000;
assign logo_start[16][37] = 9'b100000000;
assign logo_start[17][3] = 9'b100000000;
assign logo_start[17][4] = 9'b100000000;
assign logo_start[17][5] = 9'b100100000;
assign logo_start[17][6] = 9'b100100000;
assign logo_start[17][7] = 9'b100100000;
assign logo_start[17][8] = 9'b100100000;
assign logo_start[17][9] = 9'b100100000;
assign logo_start[17][10] = 9'b100100000;
assign logo_start[17][11] = 9'b100100000;
assign logo_start[17][12] = 9'b100100000;
assign logo_start[17][13] = 9'b100100000;
assign logo_start[17][14] = 9'b100100000;
assign logo_start[17][15] = 9'b100100000;
assign logo_start[17][16] = 9'b100100000;
assign logo_start[17][17] = 9'b100100000;
assign logo_start[17][18] = 9'b100100000;
assign logo_start[17][19] = 9'b100100000;
assign logo_start[17][20] = 9'b100100000;
assign logo_start[17][21] = 9'b100100000;
assign logo_start[17][22] = 9'b100100000;
assign logo_start[17][23] = 9'b100100000;
assign logo_start[17][24] = 9'b100100000;
assign logo_start[17][25] = 9'b100100000;
assign logo_start[17][26] = 9'b100100000;
assign logo_start[17][27] = 9'b100100000;
assign logo_start[17][28] = 9'b100100000;
assign logo_start[17][29] = 9'b100100000;
assign logo_start[17][30] = 9'b100100000;
assign logo_start[17][31] = 9'b100100000;
assign logo_start[17][32] = 9'b100100000;
assign logo_start[17][33] = 9'b100100000;
assign logo_start[17][34] = 9'b100100000;
assign logo_start[17][35] = 9'b100000000;
assign logo_start[17][36] = 9'b100000000;
assign logo_start[18][5] = 9'b100000000;
assign logo_start[18][6] = 9'b100000000;
assign logo_start[18][7] = 9'b100000000;
assign logo_start[18][8] = 9'b100000000;
assign logo_start[18][9] = 9'b100000000;
assign logo_start[18][10] = 9'b100000000;
assign logo_start[18][11] = 9'b100000000;
assign logo_start[18][12] = 9'b100000000;
assign logo_start[18][13] = 9'b100000000;
assign logo_start[18][14] = 9'b100000000;
assign logo_start[18][15] = 9'b100000000;
assign logo_start[18][16] = 9'b100000000;
assign logo_start[18][17] = 9'b100000000;
assign logo_start[18][18] = 9'b100000000;
assign logo_start[18][19] = 9'b100000000;
assign logo_start[18][20] = 9'b100000000;
assign logo_start[18][21] = 9'b100000000;
assign logo_start[18][22] = 9'b100000000;
assign logo_start[18][23] = 9'b100000000;
assign logo_start[18][24] = 9'b100000000;
assign logo_start[18][25] = 9'b100000000;
assign logo_start[18][26] = 9'b100000000;
assign logo_start[18][27] = 9'b100000000;
assign logo_start[18][28] = 9'b100000000;
assign logo_start[18][29] = 9'b100000000;
assign logo_start[18][30] = 9'b100000000;
assign logo_start[18][31] = 9'b100000000;
assign logo_start[18][32] = 9'b100000000;
assign logo_start[18][33] = 9'b100000000;
assign logo_start[18][34] = 9'b100000000;
assign logo_start[18][35] = 9'b100000000;
//Total de Lineas = 646
endmodule

