`timescale 1ns / 1ps
module police1 (
input enable,
input clock,
input [9:0] posx, posy,
input [9:0] hcount,
input [9:0] vcount,
output reg[2:0] red,
output reg[2:0] green,
output reg[1:0] blue,
output reg data);

always @(posedge clock)
begin
	if(enable)
	begin
		if(hcount >= posx & hcount < posx + RESOLUCION_X & vcount >= posy & vcount < posy + RESOLUCION_Y)
		begin
			if (police1[vcount - posy][hcount - posx][8] == 1'b1)
			begin
				red   <= police1[vcount- posy][hcount- posx][7:5];
				green <= police1[vcount- posy][hcount- posx][4:2];
            blue 	<= police1[vcount- posy][hcount- posx][1:0];
				data  <= 1'b1;
			end
			else
				data <= 0;
			end
		else
		data <= 0;
	end
end

parameter RESOLUCION_X = 18;
parameter RESOLUCION_Y = 45;
wire [8:0] police1[RESOLUCION_Y - 1'b1 : 0][RESOLUCION_X - 1'b1 : 0];
assign police1[1][5] = 9'b110110101;
assign police1[1][6] = 9'b110010001;
assign police1[1][7] = 9'b110010001;
assign police1[1][8] = 9'b101101101;
assign police1[1][9] = 9'b101101101;
assign police1[1][10] = 9'b110010001;
assign police1[1][11] = 9'b110010001;
assign police1[1][12] = 9'b110010001;
assign police1[2][3] = 9'b111111101;
assign police1[2][4] = 9'b111111110;
assign police1[2][5] = 9'b101101110;
assign police1[2][6] = 9'b101001001;
assign police1[2][7] = 9'b100100101;
assign police1[2][8] = 9'b100000001;
assign police1[2][9] = 9'b100000001;
assign police1[2][10] = 9'b100100101;
assign police1[2][11] = 9'b101001001;
assign police1[2][12] = 9'b101101101;
assign police1[2][13] = 9'b111111110;
assign police1[2][14] = 9'b111111111;
assign police1[3][2] = 9'b110110101;
assign police1[3][3] = 9'b111111101;
assign police1[3][4] = 9'b100100101;
assign police1[3][5] = 9'b100000001;
assign police1[3][6] = 9'b100000001;
assign police1[3][7] = 9'b100000001;
assign police1[3][8] = 9'b100000001;
assign police1[3][9] = 9'b100000001;
assign police1[3][10] = 9'b100000001;
assign police1[3][11] = 9'b100000001;
assign police1[3][12] = 9'b100000001;
assign police1[3][13] = 9'b100100101;
assign police1[3][14] = 9'b111111110;
assign police1[3][15] = 9'b110110101;
assign police1[4][1] = 9'b101101101;
assign police1[4][2] = 9'b110110101;
assign police1[4][3] = 9'b101101110;
assign police1[4][4] = 9'b100000001;
assign police1[4][5] = 9'b100000001;
assign police1[4][6] = 9'b100000001;
assign police1[4][7] = 9'b100000001;
assign police1[4][8] = 9'b100000001;
assign police1[4][9] = 9'b100000001;
assign police1[4][10] = 9'b100000001;
assign police1[4][11] = 9'b100000001;
assign police1[4][12] = 9'b100000001;
assign police1[4][13] = 9'b100000001;
assign police1[4][14] = 9'b101101110;
assign police1[4][15] = 9'b110110101;
assign police1[4][16] = 9'b110010001;
assign police1[5][1] = 9'b101101100;
assign police1[5][2] = 9'b110010001;
assign police1[5][3] = 9'b101101110;
assign police1[5][4] = 9'b100000001;
assign police1[5][5] = 9'b100000001;
assign police1[5][6] = 9'b100000001;
assign police1[5][7] = 9'b100000001;
assign police1[5][8] = 9'b100000001;
assign police1[5][9] = 9'b100000001;
assign police1[5][10] = 9'b100000001;
assign police1[5][11] = 9'b100000001;
assign police1[5][12] = 9'b100000001;
assign police1[5][13] = 9'b100000001;
assign police1[5][14] = 9'b101001001;
assign police1[5][15] = 9'b110010001;
assign police1[5][16] = 9'b101101101;
assign police1[6][1] = 9'b101101101;
assign police1[6][2] = 9'b110010010;
assign police1[6][3] = 9'b101001001;
assign police1[6][4] = 9'b100000001;
assign police1[6][5] = 9'b100000001;
assign police1[6][6] = 9'b100000001;
assign police1[6][7] = 9'b100000001;
assign police1[6][8] = 9'b100000001;
assign police1[6][9] = 9'b100000001;
assign police1[6][10] = 9'b100000001;
assign police1[6][11] = 9'b100000001;
assign police1[6][12] = 9'b100000001;
assign police1[6][13] = 9'b100000001;
assign police1[6][14] = 9'b100100101;
assign police1[6][15] = 9'b110010010;
assign police1[6][16] = 9'b101101101;
assign police1[7][1] = 9'b101101101;
assign police1[7][2] = 9'b110010001;
assign police1[7][3] = 9'b101001001;
assign police1[7][4] = 9'b100000001;
assign police1[7][5] = 9'b100000001;
assign police1[7][6] = 9'b100000001;
assign police1[7][7] = 9'b100000001;
assign police1[7][8] = 9'b100000001;
assign police1[7][9] = 9'b100000001;
assign police1[7][10] = 9'b100000001;
assign police1[7][11] = 9'b100000001;
assign police1[7][12] = 9'b100000001;
assign police1[7][13] = 9'b100000001;
assign police1[7][14] = 9'b100000001;
assign police1[7][15] = 9'b110010001;
assign police1[7][16] = 9'b101101101;
assign police1[8][1] = 9'b101101101;
assign police1[8][2] = 9'b110010001;
assign police1[8][3] = 9'b101001010;
assign police1[8][4] = 9'b100100101;
assign police1[8][5] = 9'b100000001;
assign police1[8][6] = 9'b100100101;
assign police1[8][7] = 9'b100100101;
assign police1[8][8] = 9'b100100101;
assign police1[8][9] = 9'b100100101;
assign police1[8][10] = 9'b100100101;
assign police1[8][11] = 9'b100100101;
assign police1[8][12] = 9'b100000001;
assign police1[8][13] = 9'b100000001;
assign police1[8][14] = 9'b100000001;
assign police1[8][15] = 9'b101101101;
assign police1[8][16] = 9'b101101101;
assign police1[9][1] = 9'b101101101;
assign police1[9][2] = 9'b101101101;
assign police1[9][3] = 9'b101001010;
assign police1[9][4] = 9'b100100101;
assign police1[9][5] = 9'b100000001;
assign police1[9][6] = 9'b100000001;
assign police1[9][7] = 9'b100000001;
assign police1[9][8] = 9'b100000001;
assign police1[9][9] = 9'b100000001;
assign police1[9][10] = 9'b100000001;
assign police1[9][11] = 9'b100000001;
assign police1[9][12] = 9'b100000001;
assign police1[9][13] = 9'b100000001;
assign police1[9][14] = 9'b100000001;
assign police1[9][15] = 9'b101101101;
assign police1[9][16] = 9'b101101101;
assign police1[10][1] = 9'b101101101;
assign police1[10][2] = 9'b101101101;
assign police1[10][3] = 9'b101001010;
assign police1[10][4] = 9'b100100101;
assign police1[10][5] = 9'b100000001;
assign police1[10][6] = 9'b100000001;
assign police1[10][7] = 9'b100000001;
assign police1[10][8] = 9'b100000001;
assign police1[10][9] = 9'b100000001;
assign police1[10][10] = 9'b100000001;
assign police1[10][11] = 9'b100000001;
assign police1[10][12] = 9'b100000001;
assign police1[10][13] = 9'b100000001;
assign police1[10][14] = 9'b100000001;
assign police1[10][15] = 9'b101001001;
assign police1[10][16] = 9'b101101101;
assign police1[11][1] = 9'b101101101;
assign police1[11][2] = 9'b101101110;
assign police1[11][3] = 9'b101101110;
assign police1[11][4] = 9'b101001001;
assign police1[11][5] = 9'b100100101;
assign police1[11][6] = 9'b100000001;
assign police1[11][7] = 9'b100000001;
assign police1[11][8] = 9'b100000001;
assign police1[11][9] = 9'b100000001;
assign police1[11][10] = 9'b100000001;
assign police1[11][11] = 9'b100000001;
assign police1[11][12] = 9'b100000001;
assign police1[11][13] = 9'b100000001;
assign police1[11][14] = 9'b100000001;
assign police1[11][15] = 9'b101001001;
assign police1[11][16] = 9'b101101101;
assign police1[12][1] = 9'b101101101;
assign police1[12][2] = 9'b101101110;
assign police1[12][3] = 9'b101101110;
assign police1[12][4] = 9'b101001001;
assign police1[12][5] = 9'b100100101;
assign police1[12][6] = 9'b100000001;
assign police1[12][7] = 9'b100000001;
assign police1[12][8] = 9'b100000001;
assign police1[12][9] = 9'b100000001;
assign police1[12][10] = 9'b100000001;
assign police1[12][11] = 9'b100000001;
assign police1[12][12] = 9'b100000001;
assign police1[12][13] = 9'b100000001;
assign police1[12][14] = 9'b100000001;
assign police1[12][15] = 9'b100100101;
assign police1[12][16] = 9'b101101101;
assign police1[13][1] = 9'b101101101;
assign police1[13][2] = 9'b110010010;
assign police1[13][3] = 9'b101101110;
assign police1[13][4] = 9'b101001010;
assign police1[13][5] = 9'b100100101;
assign police1[13][6] = 9'b100000001;
assign police1[13][7] = 9'b100000001;
assign police1[13][8] = 9'b100000001;
assign police1[13][9] = 9'b100000001;
assign police1[13][10] = 9'b100000001;
assign police1[13][11] = 9'b100000001;
assign police1[13][12] = 9'b100000001;
assign police1[13][13] = 9'b100000001;
assign police1[13][14] = 9'b100000001;
assign police1[13][15] = 9'b100100101;
assign police1[13][16] = 9'b101101101;
assign police1[14][1] = 9'b101101101;
assign police1[14][2] = 9'b110010010;
assign police1[14][3] = 9'b101101111;
assign police1[14][4] = 9'b101001010;
assign police1[14][5] = 9'b100100101;
assign police1[14][6] = 9'b100000001;
assign police1[14][7] = 9'b100000001;
assign police1[14][8] = 9'b100000001;
assign police1[14][9] = 9'b100000001;
assign police1[14][10] = 9'b100000001;
assign police1[14][11] = 9'b100000001;
assign police1[14][12] = 9'b100000001;
assign police1[14][13] = 9'b100000001;
assign police1[14][14] = 9'b100000001;
assign police1[14][15] = 9'b100000001;
assign police1[14][16] = 9'b101101101;
assign police1[15][1] = 9'b101101101;
assign police1[15][2] = 9'b110010010;
assign police1[15][3] = 9'b110010011;
assign police1[15][4] = 9'b101101110;
assign police1[15][5] = 9'b101001001;
assign police1[15][6] = 9'b100000001;
assign police1[15][7] = 9'b100000001;
assign police1[15][8] = 9'b100000001;
assign police1[15][9] = 9'b100000001;
assign police1[15][10] = 9'b100000001;
assign police1[15][11] = 9'b100000001;
assign police1[15][12] = 9'b100000001;
assign police1[15][13] = 9'b100000001;
assign police1[15][14] = 9'b100000001;
assign police1[15][15] = 9'b100000001;
assign police1[15][16] = 9'b101101101;
assign police1[16][1] = 9'b101001001;
assign police1[16][2] = 9'b110010010;
assign police1[16][3] = 9'b110010011;
assign police1[16][4] = 9'b101001001;
assign police1[16][5] = 9'b100100101;
assign police1[16][6] = 9'b100100101;
assign police1[16][7] = 9'b100100101;
assign police1[16][8] = 9'b100100101;
assign police1[16][9] = 9'b100100101;
assign police1[16][10] = 9'b100100101;
assign police1[16][11] = 9'b100000001;
assign police1[16][12] = 9'b100000001;
assign police1[16][13] = 9'b100000001;
assign police1[16][14] = 9'b100000001;
assign police1[16][15] = 9'b100000001;
assign police1[16][16] = 9'b101001001;
assign police1[17][1] = 9'b101001001;
assign police1[17][2] = 9'b110010010;
assign police1[17][3] = 9'b101001010;
assign police1[17][4] = 9'b100100101;
assign police1[17][5] = 9'b101001010;
assign police1[17][6] = 9'b101101111;
assign police1[17][7] = 9'b110010011;
assign police1[17][8] = 9'b110110111;
assign police1[17][9] = 9'b110110111;
assign police1[17][10] = 9'b110010011;
assign police1[17][11] = 9'b101101111;
assign police1[17][12] = 9'b101001011;
assign police1[17][13] = 9'b100100101;
assign police1[17][14] = 9'b100000001;
assign police1[17][15] = 9'b100000001;
assign police1[17][16] = 9'b101001001;
assign police1[18][1] = 9'b101001000;
assign police1[18][2] = 9'b101001001;
assign police1[18][3] = 9'b100100110;
assign police1[18][4] = 9'b101101111;
assign police1[18][5] = 9'b101101111;
assign police1[18][6] = 9'b110010011;
assign police1[18][7] = 9'b110010011;
assign police1[18][8] = 9'b110010011;
assign police1[18][9] = 9'b110110111;
assign police1[18][10] = 9'b111111111;
assign police1[18][11] = 9'b110110111;
assign police1[18][12] = 9'b110010011;
assign police1[18][13] = 9'b110010011;
assign police1[18][14] = 9'b101001010;
assign police1[18][15] = 9'b100000001;
assign police1[18][16] = 9'b101001001;
assign police1[19][1] = 9'b101001001;
assign police1[19][2] = 9'b100100101;
assign police1[19][3] = 9'b110010011;
assign police1[19][4] = 9'b110010011;
assign police1[19][5] = 9'b101101110;
assign police1[19][6] = 9'b101101111;
assign police1[19][7] = 9'b110010011;
assign police1[19][8] = 9'b110010011;
assign police1[19][9] = 9'b110010011;
assign police1[19][10] = 9'b110110111;
assign police1[19][11] = 9'b111111111;
assign police1[19][12] = 9'b111111111;
assign police1[19][13] = 9'b111111111;
assign police1[19][14] = 9'b110110111;
assign police1[19][15] = 9'b101001001;
assign police1[19][16] = 9'b100000000;
assign police1[20][1] = 9'b101001001;
assign police1[20][2] = 9'b101001001;
assign police1[20][3] = 9'b110110111;
assign police1[20][4] = 9'b110010011;
assign police1[20][5] = 9'b101110011;
assign police1[20][6] = 9'b101101111;
assign police1[20][7] = 9'b110010011;
assign police1[20][8] = 9'b110010011;
assign police1[20][9] = 9'b110010011;
assign police1[20][10] = 9'b110010011;
assign police1[20][11] = 9'b110110111;
assign police1[20][12] = 9'b111111111;
assign police1[20][13] = 9'b111111111;
assign police1[20][14] = 9'b111111111;
assign police1[20][15] = 9'b100100101;
assign police1[20][16] = 9'b100000001;
assign police1[21][1] = 9'b101001001;
assign police1[21][2] = 9'b101001001;
assign police1[21][3] = 9'b110010011;
assign police1[21][4] = 9'b110110111;
assign police1[21][5] = 9'b110010111;
assign police1[21][6] = 9'b110010011;
assign police1[21][7] = 9'b110010011;
assign police1[21][8] = 9'b101101111;
assign police1[21][9] = 9'b101101111;
assign police1[21][10] = 9'b110010011;
assign police1[21][11] = 9'b110010011;
assign police1[21][12] = 9'b110010011;
assign police1[21][13] = 9'b110010011;
assign police1[21][14] = 9'b110010011;
assign police1[21][15] = 9'b101001001;
assign police1[21][16] = 9'b100000001;
assign police1[22][0] = 9'b100000000;
assign police1[22][1] = 9'b100100100;
assign police1[22][2] = 9'b101001001;
assign police1[22][3] = 9'b101101110;
assign police1[22][4] = 9'b110110111;
assign police1[22][5] = 9'b110110111;
assign police1[22][6] = 9'b110010011;
assign police1[22][7] = 9'b101101111;
assign police1[22][8] = 9'b101101110;
assign police1[22][9] = 9'b101001010;
assign police1[22][10] = 9'b101001011;
assign police1[22][11] = 9'b100100111;
assign police1[22][12] = 9'b101001011;
assign police1[22][13] = 9'b101001011;
assign police1[22][14] = 9'b101001111;
assign police1[22][15] = 9'b101001001;
assign police1[22][16] = 9'b100000000;
assign police1[22][17] = 9'b101001001;
assign police1[23][0] = 9'b100100100;
assign police1[23][1] = 9'b101001001;
assign police1[23][2] = 9'b101001001;
assign police1[23][3] = 9'b101001001;
assign police1[23][4] = 9'b110010011;
assign police1[23][5] = 9'b110010011;
assign police1[23][6] = 9'b110010011;
assign police1[23][7] = 9'b110010011;
assign police1[23][8] = 9'b101101111;
assign police1[23][9] = 9'b101101110;
assign police1[23][10] = 9'b101001010;
assign police1[23][11] = 9'b101001010;
assign police1[23][12] = 9'b100100110;
assign police1[23][13] = 9'b100100111;
assign police1[23][14] = 9'b101001010;
assign police1[23][15] = 9'b101001001;
assign police1[23][16] = 9'b100000001;
assign police1[23][17] = 9'b101001001;
assign police1[24][1] = 9'b101001001;
assign police1[24][2] = 9'b101101101;
assign police1[24][3] = 9'b101001001;
assign police1[24][4] = 9'b101101101;
assign police1[24][5] = 9'b101101101;
assign police1[24][6] = 9'b110010001;
assign police1[24][7] = 9'b110010001;
assign police1[24][8] = 9'b110010001;
assign police1[24][9] = 9'b110010001;
assign police1[24][10] = 9'b110010001;
assign police1[24][11] = 9'b110010001;
assign police1[24][12] = 9'b101101101;
assign police1[24][13] = 9'b101101101;
assign police1[24][14] = 9'b101001001;
assign police1[24][15] = 9'b101001001;
assign police1[24][16] = 9'b100000001;
assign police1[25][1] = 9'b101001001;
assign police1[25][2] = 9'b101001001;
assign police1[25][3] = 9'b110010001;
assign police1[25][4] = 9'b110110110;
assign police1[25][5] = 9'b110010010;
assign police1[25][6] = 9'b110010010;
assign police1[25][7] = 9'b110010010;
assign police1[25][8] = 9'b110010010;
assign police1[25][9] = 9'b110010010;
assign police1[25][10] = 9'b110010010;
assign police1[25][11] = 9'b110010010;
assign police1[25][12] = 9'b110110110;
assign police1[25][13] = 9'b110110110;
assign police1[25][14] = 9'b101101101;
assign police1[25][15] = 9'b101001001;
assign police1[25][16] = 9'b100000001;
assign police1[26][1] = 9'b101001001;
assign police1[26][2] = 9'b101001001;
assign police1[26][3] = 9'b101101101;
assign police1[26][4] = 9'b110010001;
assign police1[26][5] = 9'b110010001;
assign police1[26][6] = 9'b110010001;
assign police1[26][7] = 9'b110010001;
assign police1[26][8] = 9'b110010001;
assign police1[26][9] = 9'b110010001;
assign police1[26][10] = 9'b110010001;
assign police1[26][11] = 9'b110010001;
assign police1[26][12] = 9'b110010001;
assign police1[26][13] = 9'b110010010;
assign police1[26][14] = 9'b101101101;
assign police1[26][15] = 9'b101001001;
assign police1[26][16] = 9'b100000001;
assign police1[27][1] = 9'b101001001;
assign police1[27][2] = 9'b101101101;
assign police1[27][3] = 9'b101101101;
assign police1[27][4] = 9'b110010001;
assign police1[27][5] = 9'b110010001;
assign police1[27][6] = 9'b110010001;
assign police1[27][7] = 9'b101110001;
assign police1[27][8] = 9'b101101101;
assign police1[27][9] = 9'b101101101;
assign police1[27][10] = 9'b101101101;
assign police1[27][11] = 9'b101101101;
assign police1[27][12] = 9'b110010001;
assign police1[27][13] = 9'b110010001;
assign police1[27][14] = 9'b101001001;
assign police1[27][15] = 9'b101001001;
assign police1[27][16] = 9'b100000001;
assign police1[28][1] = 9'b101001001;
assign police1[28][2] = 9'b101101101;
assign police1[28][3] = 9'b101101001;
assign police1[28][4] = 9'b101101101;
assign police1[28][5] = 9'b101001110;
assign police1[28][6] = 9'b101101001;
assign police1[28][7] = 9'b110001001;
assign police1[28][8] = 9'b110010001;
assign police1[28][9] = 9'b110010010;
assign police1[28][10] = 9'b110010010;
assign police1[28][11] = 9'b110010010;
assign police1[28][12] = 9'b101001110;
assign police1[28][13] = 9'b101101101;
assign police1[28][14] = 9'b101001001;
assign police1[28][15] = 9'b101001001;
assign police1[28][16] = 9'b100000001;
assign police1[29][1] = 9'b101001001;
assign police1[29][2] = 9'b101101101;
assign police1[29][3] = 9'b101101101;
assign police1[29][4] = 9'b101001101;
assign police1[29][5] = 9'b100001011;
assign police1[29][6] = 9'b110000000;
assign police1[29][7] = 9'b111100000;
assign police1[29][8] = 9'b111110001;
assign police1[29][9] = 9'b111111111;
assign police1[29][10] = 9'b111111111;
assign police1[29][11] = 9'b110010111;
assign police1[29][12] = 9'b100000111;
assign police1[29][13] = 9'b100101010;
assign police1[29][14] = 9'b101101101;
assign police1[29][15] = 9'b101001001;
assign police1[29][16] = 9'b100000001;
assign police1[30][1] = 9'b101101101;
assign police1[30][2] = 9'b101101101;
assign police1[30][3] = 9'b101001001;
assign police1[30][4] = 9'b101001001;
assign police1[30][5] = 9'b100000011;
assign police1[30][6] = 9'b101100000;
assign police1[30][7] = 9'b110100000;
assign police1[30][8] = 9'b110001101;
assign police1[30][9] = 9'b110010110;
assign police1[30][10] = 9'b110110110;
assign police1[30][11] = 9'b101101110;
assign police1[30][12] = 9'b100000010;
assign police1[30][13] = 9'b100101001;
assign police1[30][14] = 9'b101101101;
assign police1[30][15] = 9'b101001001;
assign police1[30][16] = 9'b100100101;
assign police1[31][1] = 9'b110010010;
assign police1[31][2] = 9'b101101101;
assign police1[31][3] = 9'b101001001;
assign police1[31][4] = 9'b101001001;
assign police1[31][5] = 9'b101001001;
assign police1[31][6] = 9'b101001001;
assign police1[31][7] = 9'b101001001;
assign police1[31][8] = 9'b101001001;
assign police1[31][9] = 9'b101001001;
assign police1[31][10] = 9'b101001001;
assign police1[31][11] = 9'b101001001;
assign police1[31][12] = 9'b101001001;
assign police1[31][13] = 9'b101001001;
assign police1[31][14] = 9'b101001001;
assign police1[31][15] = 9'b101101101;
assign police1[31][16] = 9'b100100100;
assign police1[32][1] = 9'b110010001;
assign police1[32][2] = 9'b101101101;
assign police1[32][3] = 9'b101001001;
assign police1[32][4] = 9'b100100100;
assign police1[32][5] = 9'b101001000;
assign police1[32][6] = 9'b101001000;
assign police1[32][7] = 9'b101001000;
assign police1[32][8] = 9'b101001000;
assign police1[32][9] = 9'b101001000;
assign police1[32][10] = 9'b101001000;
assign police1[32][11] = 9'b101001000;
assign police1[32][12] = 9'b101001000;
assign police1[32][13] = 9'b101001000;
assign police1[32][14] = 9'b101001001;
assign police1[32][15] = 9'b101101101;
assign police1[32][16] = 9'b101001001;
assign police1[33][1] = 9'b110010010;
assign police1[33][2] = 9'b101001001;
assign police1[33][3] = 9'b101001001;
assign police1[33][4] = 9'b101001001;
assign police1[33][5] = 9'b101001001;
assign police1[33][6] = 9'b101001001;
assign police1[33][7] = 9'b101001001;
assign police1[33][8] = 9'b101001001;
assign police1[33][9] = 9'b101001001;
assign police1[33][10] = 9'b101001001;
assign police1[33][11] = 9'b101001001;
assign police1[33][12] = 9'b101001001;
assign police1[33][13] = 9'b101001000;
assign police1[33][14] = 9'b101000100;
assign police1[33][15] = 9'b101001001;
assign police1[33][16] = 9'b101101101;
assign police1[34][1] = 9'b110010010;
assign police1[34][2] = 9'b101101101;
assign police1[34][3] = 9'b101001001;
assign police1[34][4] = 9'b110010011;
assign police1[34][5] = 9'b110010011;
assign police1[34][6] = 9'b110110111;
assign police1[34][7] = 9'b110110111;
assign police1[34][8] = 9'b110010011;
assign police1[34][9] = 9'b110010011;
assign police1[34][10] = 9'b110010011;
assign police1[34][11] = 9'b110010011;
assign police1[34][12] = 9'b110010010;
assign police1[34][13] = 9'b110010011;
assign police1[34][14] = 9'b101101101;
assign police1[34][15] = 9'b101001000;
assign police1[34][16] = 9'b101101101;
assign police1[35][1] = 9'b110010001;
assign police1[35][2] = 9'b110110110;
assign police1[35][3] = 9'b101001001;
assign police1[35][4] = 9'b101001010;
assign police1[35][5] = 9'b101101110;
assign police1[35][6] = 9'b101101110;
assign police1[35][7] = 9'b110010010;
assign police1[35][8] = 9'b110010010;
assign police1[35][9] = 9'b110010011;
assign police1[35][10] = 9'b110010011;
assign police1[35][11] = 9'b110010011;
assign police1[35][12] = 9'b110010011;
assign police1[35][13] = 9'b110010011;
assign police1[35][14] = 9'b110010010;
assign police1[35][15] = 9'b101101101;
assign police1[35][16] = 9'b101101101;
assign police1[36][1] = 9'b110010001;
assign police1[36][2] = 9'b110110111;
assign police1[36][3] = 9'b101101110;
assign police1[36][4] = 9'b101101101;
assign police1[36][5] = 9'b101101101;
assign police1[36][6] = 9'b101101110;
assign police1[36][7] = 9'b101101110;
assign police1[36][8] = 9'b101101110;
assign police1[36][9] = 9'b101101110;
assign police1[36][10] = 9'b110010010;
assign police1[36][11] = 9'b110010010;
assign police1[36][12] = 9'b110010010;
assign police1[36][13] = 9'b101101101;
assign police1[36][14] = 9'b101001001;
assign police1[36][15] = 9'b101101101;
assign police1[36][16] = 9'b101101101;
assign police1[37][1] = 9'b110010001;
assign police1[37][2] = 9'b110010010;
assign police1[37][3] = 9'b100000001;
assign police1[37][4] = 9'b100100101;
assign police1[37][5] = 9'b100100101;
assign police1[37][6] = 9'b100100101;
assign police1[37][7] = 9'b100100101;
assign police1[37][8] = 9'b100100101;
assign police1[37][9] = 9'b100100101;
assign police1[37][10] = 9'b100100101;
assign police1[37][11] = 9'b100100101;
assign police1[37][12] = 9'b100100101;
assign police1[37][13] = 9'b100000001;
assign police1[37][14] = 9'b100000001;
assign police1[37][15] = 9'b101001001;
assign police1[37][16] = 9'b101101101;
assign police1[38][1] = 9'b101101101;
assign police1[38][2] = 9'b110010010;
assign police1[38][3] = 9'b100000001;
assign police1[38][4] = 9'b100000001;
assign police1[38][5] = 9'b100000001;
assign police1[38][6] = 9'b100000001;
assign police1[38][7] = 9'b100000001;
assign police1[38][8] = 9'b100000001;
assign police1[38][9] = 9'b100000001;
assign police1[38][10] = 9'b100000001;
assign police1[38][11] = 9'b100000001;
assign police1[38][12] = 9'b100000001;
assign police1[38][13] = 9'b100000001;
assign police1[38][14] = 9'b100000001;
assign police1[38][15] = 9'b101101101;
assign police1[38][16] = 9'b101101101;
assign police1[39][1] = 9'b101101101;
assign police1[39][2] = 9'b110110110;
assign police1[39][3] = 9'b100100101;
assign police1[39][4] = 9'b100000001;
assign police1[39][5] = 9'b100000001;
assign police1[39][6] = 9'b100000001;
assign police1[39][7] = 9'b100000001;
assign police1[39][8] = 9'b100000001;
assign police1[39][9] = 9'b100000001;
assign police1[39][10] = 9'b100000001;
assign police1[39][11] = 9'b100000001;
assign police1[39][12] = 9'b100000001;
assign police1[39][13] = 9'b100000001;
assign police1[39][14] = 9'b100000001;
assign police1[39][15] = 9'b101101101;
assign police1[39][16] = 9'b101101101;
assign police1[40][1] = 9'b101101101;
assign police1[40][2] = 9'b110110110;
assign police1[40][3] = 9'b101101110;
assign police1[40][4] = 9'b100000001;
assign police1[40][5] = 9'b100000001;
assign police1[40][6] = 9'b100000001;
assign police1[40][7] = 9'b100000001;
assign police1[40][8] = 9'b100000001;
assign police1[40][9] = 9'b100000001;
assign police1[40][10] = 9'b100000001;
assign police1[40][11] = 9'b100000001;
assign police1[40][12] = 9'b100000001;
assign police1[40][13] = 9'b100000001;
assign police1[40][14] = 9'b100100101;
assign police1[40][15] = 9'b101101101;
assign police1[40][16] = 9'b101101101;
assign police1[41][2] = 9'b110010001;
assign police1[41][3] = 9'b110110010;
assign police1[41][4] = 9'b100000001;
assign police1[41][5] = 9'b100000001;
assign police1[41][6] = 9'b100000001;
assign police1[41][7] = 9'b100000001;
assign police1[41][8] = 9'b100000001;
assign police1[41][9] = 9'b100000001;
assign police1[41][10] = 9'b100000001;
assign police1[41][11] = 9'b100000001;
assign police1[41][12] = 9'b100000001;
assign police1[41][13] = 9'b100000001;
assign police1[41][14] = 9'b110001101;
assign police1[41][15] = 9'b110001101;
assign police1[42][3] = 9'b111110110;
assign police1[42][4] = 9'b110110110;
assign police1[42][5] = 9'b101101110;
assign police1[42][6] = 9'b101001010;
assign police1[42][7] = 9'b101001001;
assign police1[42][8] = 9'b100100101;
assign police1[42][9] = 9'b100100101;
assign police1[42][10] = 9'b101001001;
assign police1[42][11] = 9'b101001010;
assign police1[42][12] = 9'b101101110;
assign police1[42][13] = 9'b110010010;
assign police1[42][14] = 9'b111110110;
assign police1[43][5] = 9'b111111111;
assign police1[43][6] = 9'b111111111;
assign police1[43][7] = 9'b111111111;
assign police1[43][8] = 9'b111111111;
assign police1[43][9] = 9'b111111111;
assign police1[43][10] = 9'b111111111;
assign police1[43][11] = 9'b111111111;
assign police1[43][12] = 9'b111111111;
//Total de Lineas = 664
endmodule

