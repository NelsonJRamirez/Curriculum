`timescale 1ns / 1ps
module ferrary (
input enable,
input clock,
input [9:0] posx, posy,
input [9:0] hcount,
input [9:0] vcount,
output reg[2:0] red,
output reg[2:0] green,
output reg[1:0] blue,
output reg data);

always @(posedge clock)
begin
	if(enable)
	begin
		if(hcount >= posx & hcount < posx + RESOLUCION_X & vcount >= posy & vcount < posy + RESOLUCION_Y)
		begin
			if (ferrary[vcount - posy][hcount - posx][8] == 1'b1)
			begin
				red   <= ferrary[vcount- posy][hcount- posx][7:5];
				green <= ferrary[vcount- posy][hcount- posx][4:2];
            blue 	<= ferrary[vcount- posy][hcount- posx][1:0];
				data  <= 1'b1;
			end
			else
				data <= 0;
			end
		else
		data <= 0;
	end
end

parameter RESOLUCION_X = 25;
parameter RESOLUCION_Y = 50;
wire [8:0] ferrary[RESOLUCION_Y - 1'b1 : 0][RESOLUCION_X - 1'b1 : 0];
assign ferrary[3][8] = 9'b100000000;
assign ferrary[3][9] = 9'b100000000;
assign ferrary[3][10] = 9'b100000100;
assign ferrary[3][11] = 9'b100100101;
assign ferrary[3][12] = 9'b100100101;
assign ferrary[3][13] = 9'b100000100;
assign ferrary[3][14] = 9'b100000100;
assign ferrary[3][15] = 9'b100000000;
assign ferrary[4][6] = 9'b100000000;
assign ferrary[4][7] = 9'b100100100;
assign ferrary[4][8] = 9'b100101001;
assign ferrary[4][9] = 9'b100101001;
assign ferrary[4][10] = 9'b101001101;
assign ferrary[4][11] = 9'b101001101;
assign ferrary[4][12] = 9'b101101110;
assign ferrary[4][13] = 9'b101001110;
assign ferrary[4][14] = 9'b101001101;
assign ferrary[4][15] = 9'b101001001;
assign ferrary[4][16] = 9'b100100100;
assign ferrary[4][17] = 9'b100100000;
assign ferrary[5][5] = 9'b100100100;
assign ferrary[5][6] = 9'b100100000;
assign ferrary[5][7] = 9'b101001001;
assign ferrary[5][8] = 9'b101001001;
assign ferrary[5][9] = 9'b101001101;
assign ferrary[5][10] = 9'b101001110;
assign ferrary[5][11] = 9'b101101110;
assign ferrary[5][12] = 9'b101110010;
assign ferrary[5][13] = 9'b101101110;
assign ferrary[5][14] = 9'b101001110;
assign ferrary[5][15] = 9'b101001110;
assign ferrary[5][16] = 9'b101001001;
assign ferrary[5][17] = 9'b101000000;
assign ferrary[5][18] = 9'b100100101;
assign ferrary[6][4] = 9'b100000000;
assign ferrary[6][5] = 9'b100100100;
assign ferrary[6][6] = 9'b100100000;
assign ferrary[6][7] = 9'b100101001;
assign ferrary[6][8] = 9'b100101001;
assign ferrary[6][9] = 9'b101001001;
assign ferrary[6][10] = 9'b101001101;
assign ferrary[6][11] = 9'b101001101;
assign ferrary[6][12] = 9'b101001101;
assign ferrary[6][13] = 9'b101001101;
assign ferrary[6][14] = 9'b101001101;
assign ferrary[6][15] = 9'b101001101;
assign ferrary[6][16] = 9'b101001001;
assign ferrary[6][17] = 9'b101000100;
assign ferrary[6][18] = 9'b101001001;
assign ferrary[6][19] = 9'b100000000;
assign ferrary[7][4] = 9'b100100100;
assign ferrary[7][5] = 9'b100101001;
assign ferrary[7][6] = 9'b100100101;
assign ferrary[7][7] = 9'b100101001;
assign ferrary[7][8] = 9'b100101001;
assign ferrary[7][9] = 9'b100101001;
assign ferrary[7][10] = 9'b100101001;
assign ferrary[7][11] = 9'b100101001;
assign ferrary[7][12] = 9'b101001001;
assign ferrary[7][13] = 9'b101001001;
assign ferrary[7][14] = 9'b101001001;
assign ferrary[7][15] = 9'b100101001;
assign ferrary[7][16] = 9'b101001001;
assign ferrary[7][17] = 9'b101001001;
assign ferrary[7][18] = 9'b101101110;
assign ferrary[7][19] = 9'b100100101;
assign ferrary[8][4] = 9'b100101001;
assign ferrary[8][5] = 9'b101001001;
assign ferrary[8][6] = 9'b101001001;
assign ferrary[8][7] = 9'b100101001;
assign ferrary[8][8] = 9'b100100101;
assign ferrary[8][9] = 9'b100100101;
assign ferrary[8][10] = 9'b100101001;
assign ferrary[8][11] = 9'b100101001;
assign ferrary[8][12] = 9'b100101001;
assign ferrary[8][13] = 9'b100101001;
assign ferrary[8][14] = 9'b100101001;
assign ferrary[8][15] = 9'b100101001;
assign ferrary[8][16] = 9'b100101001;
assign ferrary[8][17] = 9'b101001101;
assign ferrary[8][18] = 9'b110010011;
assign ferrary[8][19] = 9'b101001001;
assign ferrary[9][4] = 9'b101001001;
assign ferrary[9][5] = 9'b101001001;
assign ferrary[9][6] = 9'b101001101;
assign ferrary[9][7] = 9'b100100101;
assign ferrary[9][8] = 9'b100100101;
assign ferrary[9][9] = 9'b100100101;
assign ferrary[9][10] = 9'b100100101;
assign ferrary[9][11] = 9'b100100101;
assign ferrary[9][12] = 9'b100100101;
assign ferrary[9][13] = 9'b100100101;
assign ferrary[9][14] = 9'b100100101;
assign ferrary[9][15] = 9'b100100101;
assign ferrary[9][16] = 9'b100100101;
assign ferrary[9][17] = 9'b101001101;
assign ferrary[9][18] = 9'b110010111;
assign ferrary[9][19] = 9'b101101101;
assign ferrary[10][4] = 9'b101001101;
assign ferrary[10][5] = 9'b101001101;
assign ferrary[10][6] = 9'b101001101;
assign ferrary[10][7] = 9'b100100101;
assign ferrary[10][8] = 9'b100100101;
assign ferrary[10][9] = 9'b100101001;
assign ferrary[10][10] = 9'b100101001;
assign ferrary[10][11] = 9'b101001001;
assign ferrary[10][12] = 9'b100101001;
assign ferrary[10][13] = 9'b100101001;
assign ferrary[10][14] = 9'b100100101;
assign ferrary[10][15] = 9'b100100101;
assign ferrary[10][16] = 9'b100100101;
assign ferrary[10][17] = 9'b101001001;
assign ferrary[10][18] = 9'b110010111;
assign ferrary[10][19] = 9'b110010010;
assign ferrary[11][4] = 9'b101101101;
assign ferrary[11][5] = 9'b101110010;
assign ferrary[11][6] = 9'b101101110;
assign ferrary[11][7] = 9'b100101001;
assign ferrary[11][8] = 9'b100101001;
assign ferrary[11][9] = 9'b100101001;
assign ferrary[11][10] = 9'b100101001;
assign ferrary[11][11] = 9'b100101001;
assign ferrary[11][12] = 9'b100101001;
assign ferrary[11][13] = 9'b100101001;
assign ferrary[11][14] = 9'b100100101;
assign ferrary[11][15] = 9'b100100101;
assign ferrary[11][16] = 9'b100101001;
assign ferrary[11][17] = 9'b101001001;
assign ferrary[11][18] = 9'b110010111;
assign ferrary[11][19] = 9'b110111111;
assign ferrary[11][20] = 9'b100100100;
assign ferrary[12][3] = 9'b100000000;
assign ferrary[12][4] = 9'b101101101;
assign ferrary[12][5] = 9'b110010111;
assign ferrary[12][6] = 9'b101001101;
assign ferrary[12][7] = 9'b100100101;
assign ferrary[12][8] = 9'b100100101;
assign ferrary[12][9] = 9'b100100101;
assign ferrary[12][10] = 9'b100100101;
assign ferrary[12][11] = 9'b100100101;
assign ferrary[12][12] = 9'b100100101;
assign ferrary[12][13] = 9'b100100101;
assign ferrary[12][14] = 9'b100100101;
assign ferrary[12][15] = 9'b100100101;
assign ferrary[12][16] = 9'b100101001;
assign ferrary[12][17] = 9'b100101001;
assign ferrary[12][18] = 9'b110010010;
assign ferrary[12][19] = 9'b111111111;
assign ferrary[12][20] = 9'b100100100;
assign ferrary[13][3] = 9'b100000000;
assign ferrary[13][4] = 9'b101101101;
assign ferrary[13][5] = 9'b110010010;
assign ferrary[13][6] = 9'b101001001;
assign ferrary[13][7] = 9'b100101001;
assign ferrary[13][8] = 9'b101001001;
assign ferrary[13][9] = 9'b101001001;
assign ferrary[13][10] = 9'b101001101;
assign ferrary[13][11] = 9'b101101101;
assign ferrary[13][12] = 9'b101101101;
assign ferrary[13][13] = 9'b101001101;
assign ferrary[13][14] = 9'b101101101;
assign ferrary[13][15] = 9'b101001101;
assign ferrary[13][16] = 9'b101001001;
assign ferrary[13][17] = 9'b101001001;
assign ferrary[13][18] = 9'b110010010;
assign ferrary[13][19] = 9'b111111111;
assign ferrary[13][20] = 9'b100100100;
assign ferrary[14][4] = 9'b101001001;
assign ferrary[14][5] = 9'b101101101;
assign ferrary[14][6] = 9'b110001101;
assign ferrary[14][7] = 9'b110110101;
assign ferrary[14][8] = 9'b110110001;
assign ferrary[14][9] = 9'b111110101;
assign ferrary[14][10] = 9'b111110101;
assign ferrary[14][11] = 9'b111110110;
assign ferrary[14][12] = 9'b111111110;
assign ferrary[14][13] = 9'b111110101;
assign ferrary[14][14] = 9'b110010001;
assign ferrary[14][15] = 9'b110010001;
assign ferrary[14][16] = 9'b111110101;
assign ferrary[14][17] = 9'b110001101;
assign ferrary[14][18] = 9'b101101101;
assign ferrary[14][19] = 9'b110111111;
assign ferrary[14][20] = 9'b100100100;
assign ferrary[15][4] = 9'b100101001;
assign ferrary[15][5] = 9'b101101101;
assign ferrary[15][6] = 9'b110110001;
assign ferrary[15][7] = 9'b110010001;
assign ferrary[15][8] = 9'b110001101;
assign ferrary[15][9] = 9'b110001101;
assign ferrary[15][10] = 9'b110001101;
assign ferrary[15][11] = 9'b110010001;
assign ferrary[15][12] = 9'b110110001;
assign ferrary[15][13] = 9'b110001101;
assign ferrary[15][14] = 9'b101101000;
assign ferrary[15][15] = 9'b101001000;
assign ferrary[15][16] = 9'b110010001;
assign ferrary[15][17] = 9'b111111110;
assign ferrary[15][18] = 9'b101101101;
assign ferrary[15][19] = 9'b110010011;
assign ferrary[16][4] = 9'b100101001;
assign ferrary[16][5] = 9'b101001001;
assign ferrary[16][6] = 9'b110110001;
assign ferrary[16][7] = 9'b110010001;
assign ferrary[16][8] = 9'b110010001;
assign ferrary[16][9] = 9'b110010001;
assign ferrary[16][10] = 9'b101001000;
assign ferrary[16][11] = 9'b110010001;
assign ferrary[16][12] = 9'b110010001;
assign ferrary[16][13] = 9'b101001000;
assign ferrary[16][14] = 9'b101101000;
assign ferrary[16][15] = 9'b101001000;
assign ferrary[16][16] = 9'b101101000;
assign ferrary[16][17] = 9'b111111110;
assign ferrary[16][18] = 9'b101110001;
assign ferrary[16][19] = 9'b101001101;
assign ferrary[17][4] = 9'b100100101;
assign ferrary[17][5] = 9'b101001001;
assign ferrary[17][6] = 9'b110110001;
assign ferrary[17][7] = 9'b110010001;
assign ferrary[17][8] = 9'b110001101;
assign ferrary[17][9] = 9'b110010001;
assign ferrary[17][10] = 9'b101001000;
assign ferrary[17][11] = 9'b110001101;
assign ferrary[17][12] = 9'b110010001;
assign ferrary[17][13] = 9'b101001000;
assign ferrary[17][14] = 9'b101101100;
assign ferrary[17][15] = 9'b101001000;
assign ferrary[17][16] = 9'b101001000;
assign ferrary[17][17] = 9'b111111110;
assign ferrary[17][18] = 9'b110010001;
assign ferrary[17][19] = 9'b101001001;
assign ferrary[18][4] = 9'b100101001;
assign ferrary[18][5] = 9'b101001001;
assign ferrary[18][6] = 9'b110110001;
assign ferrary[18][7] = 9'b110010001;
assign ferrary[18][8] = 9'b110010001;
assign ferrary[18][9] = 9'b110110001;
assign ferrary[18][10] = 9'b110001101;
assign ferrary[18][11] = 9'b110001101;
assign ferrary[18][12] = 9'b110110001;
assign ferrary[18][13] = 9'b101101101;
assign ferrary[18][14] = 9'b101101100;
assign ferrary[18][15] = 9'b101101100;
assign ferrary[18][16] = 9'b101101000;
assign ferrary[18][17] = 9'b110010001;
assign ferrary[18][18] = 9'b110001101;
assign ferrary[18][19] = 9'b101001001;
assign ferrary[19][4] = 9'b101001001;
assign ferrary[19][5] = 9'b101001001;
assign ferrary[19][6] = 9'b110001101;
assign ferrary[19][7] = 9'b101101100;
assign ferrary[19][8] = 9'b110001101;
assign ferrary[19][9] = 9'b110001101;
assign ferrary[19][10] = 9'b101101101;
assign ferrary[19][11] = 9'b110001101;
assign ferrary[19][12] = 9'b110010001;
assign ferrary[19][13] = 9'b101101100;
assign ferrary[19][14] = 9'b101101100;
assign ferrary[19][15] = 9'b101101101;
assign ferrary[19][16] = 9'b101001000;
assign ferrary[19][17] = 9'b101101101;
assign ferrary[19][18] = 9'b101101101;
assign ferrary[19][19] = 9'b101001101;
assign ferrary[20][4] = 9'b101001001;
assign ferrary[20][5] = 9'b101101101;
assign ferrary[20][6] = 9'b101101101;
assign ferrary[20][7] = 9'b101101000;
assign ferrary[20][8] = 9'b110010001;
assign ferrary[20][9] = 9'b110010001;
assign ferrary[20][10] = 9'b101001000;
assign ferrary[20][11] = 9'b101101101;
assign ferrary[20][12] = 9'b110001101;
assign ferrary[20][13] = 9'b101000100;
assign ferrary[20][14] = 9'b110010001;
assign ferrary[20][15] = 9'b110010001;
assign ferrary[20][16] = 9'b101101101;
assign ferrary[20][17] = 9'b101101000;
assign ferrary[20][18] = 9'b110010001;
assign ferrary[20][19] = 9'b101001101;
assign ferrary[21][4] = 9'b100100101;
assign ferrary[21][5] = 9'b101101101;
assign ferrary[21][6] = 9'b101101101;
assign ferrary[21][7] = 9'b101101101;
assign ferrary[21][8] = 9'b110110001;
assign ferrary[21][9] = 9'b110110101;
assign ferrary[21][10] = 9'b101101101;
assign ferrary[21][11] = 9'b101101000;
assign ferrary[21][12] = 9'b101101101;
assign ferrary[21][13] = 9'b101101000;
assign ferrary[21][14] = 9'b110110001;
assign ferrary[21][15] = 9'b110010001;
assign ferrary[21][16] = 9'b110010001;
assign ferrary[21][17] = 9'b101101101;
assign ferrary[21][18] = 9'b110010001;
assign ferrary[21][19] = 9'b101001001;
assign ferrary[22][4] = 9'b100100100;
assign ferrary[22][5] = 9'b101101101;
assign ferrary[22][6] = 9'b101101101;
assign ferrary[22][7] = 9'b110001101;
assign ferrary[22][8] = 9'b110110101;
assign ferrary[22][9] = 9'b111111110;
assign ferrary[22][10] = 9'b110010001;
assign ferrary[22][11] = 9'b101101101;
assign ferrary[22][12] = 9'b110001101;
assign ferrary[22][13] = 9'b110010001;
assign ferrary[22][14] = 9'b111111110;
assign ferrary[22][15] = 9'b111110110;
assign ferrary[22][16] = 9'b111110110;
assign ferrary[22][17] = 9'b101101101;
assign ferrary[22][18] = 9'b110010001;
assign ferrary[22][19] = 9'b101001001;
assign ferrary[23][4] = 9'b100100100;
assign ferrary[23][5] = 9'b101101101;
assign ferrary[23][6] = 9'b101101101;
assign ferrary[23][7] = 9'b101101000;
assign ferrary[23][8] = 9'b110001101;
assign ferrary[23][9] = 9'b110010001;
assign ferrary[23][10] = 9'b110001101;
assign ferrary[23][11] = 9'b110010001;
assign ferrary[23][12] = 9'b110110101;
assign ferrary[23][13] = 9'b110010001;
assign ferrary[23][14] = 9'b101101101;
assign ferrary[23][15] = 9'b101101100;
assign ferrary[23][16] = 9'b110001101;
assign ferrary[23][17] = 9'b101101101;
assign ferrary[23][18] = 9'b110001101;
assign ferrary[23][19] = 9'b100100100;
assign ferrary[24][4] = 9'b100100101;
assign ferrary[24][5] = 9'b101101101;
assign ferrary[24][6] = 9'b101101000;
assign ferrary[24][7] = 9'b101001000;
assign ferrary[24][8] = 9'b110001101;
assign ferrary[24][9] = 9'b110010001;
assign ferrary[24][10] = 9'b101101101;
assign ferrary[24][11] = 9'b110001101;
assign ferrary[24][12] = 9'b110001101;
assign ferrary[24][13] = 9'b101101001;
assign ferrary[24][14] = 9'b101001000;
assign ferrary[24][15] = 9'b100100000;
assign ferrary[24][16] = 9'b101000100;
assign ferrary[24][17] = 9'b101101000;
assign ferrary[24][18] = 9'b101101101;
assign ferrary[24][19] = 9'b100100100;
assign ferrary[25][4] = 9'b100100101;
assign ferrary[25][5] = 9'b101101101;
assign ferrary[25][6] = 9'b100100100;
assign ferrary[25][7] = 9'b100000000;
assign ferrary[25][8] = 9'b100000000;
assign ferrary[25][9] = 9'b100000000;
assign ferrary[25][10] = 9'b100000000;
assign ferrary[25][11] = 9'b100000000;
assign ferrary[25][12] = 9'b100000000;
assign ferrary[25][13] = 9'b100100000;
assign ferrary[25][14] = 9'b100000000;
assign ferrary[25][15] = 9'b100000000;
assign ferrary[25][16] = 9'b100000000;
assign ferrary[25][17] = 9'b100100100;
assign ferrary[25][18] = 9'b101101101;
assign ferrary[25][19] = 9'b100100100;
assign ferrary[26][4] = 9'b100100100;
assign ferrary[26][5] = 9'b101101101;
assign ferrary[26][6] = 9'b100100100;
assign ferrary[26][7] = 9'b100000000;
assign ferrary[26][8] = 9'b100100000;
assign ferrary[26][9] = 9'b100100100;
assign ferrary[26][10] = 9'b100000000;
assign ferrary[26][11] = 9'b100000000;
assign ferrary[26][12] = 9'b100000000;
assign ferrary[26][13] = 9'b100000000;
assign ferrary[26][14] = 9'b100000000;
assign ferrary[26][15] = 9'b100000000;
assign ferrary[26][16] = 9'b100000000;
assign ferrary[26][17] = 9'b100100100;
assign ferrary[26][18] = 9'b101101101;
assign ferrary[26][19] = 9'b100100100;
assign ferrary[27][3] = 9'b100100101;
assign ferrary[27][4] = 9'b100100100;
assign ferrary[27][5] = 9'b101001001;
assign ferrary[27][6] = 9'b100000000;
assign ferrary[27][7] = 9'b100100100;
assign ferrary[27][8] = 9'b101001000;
assign ferrary[27][9] = 9'b101101101;
assign ferrary[27][10] = 9'b101001000;
assign ferrary[27][11] = 9'b100000000;
assign ferrary[27][12] = 9'b100000000;
assign ferrary[27][13] = 9'b101001000;
assign ferrary[27][14] = 9'b101000100;
assign ferrary[27][15] = 9'b101001000;
assign ferrary[27][16] = 9'b101000100;
assign ferrary[27][17] = 9'b101001001;
assign ferrary[27][18] = 9'b101001001;
assign ferrary[27][19] = 9'b100100100;
assign ferrary[27][20] = 9'b100101001;
assign ferrary[28][3] = 9'b100101001;
assign ferrary[28][4] = 9'b101101101;
assign ferrary[28][5] = 9'b100101001;
assign ferrary[28][6] = 9'b100100100;
assign ferrary[28][7] = 9'b100100100;
assign ferrary[28][8] = 9'b100100100;
assign ferrary[28][9] = 9'b100100100;
assign ferrary[28][10] = 9'b100100100;
assign ferrary[28][11] = 9'b100100100;
assign ferrary[28][12] = 9'b100100100;
assign ferrary[28][13] = 9'b101101000;
assign ferrary[28][14] = 9'b101000100;
assign ferrary[28][15] = 9'b100100000;
assign ferrary[28][16] = 9'b101101000;
assign ferrary[28][17] = 9'b110010001;
assign ferrary[28][18] = 9'b100101001;
assign ferrary[28][19] = 9'b101001101;
assign ferrary[28][20] = 9'b101101101;
assign ferrary[29][4] = 9'b100100101;
assign ferrary[29][5] = 9'b100101001;
assign ferrary[29][6] = 9'b101101101;
assign ferrary[29][7] = 9'b100100100;
assign ferrary[29][8] = 9'b100100100;
assign ferrary[29][9] = 9'b100100100;
assign ferrary[29][10] = 9'b100100100;
assign ferrary[29][11] = 9'b100100100;
assign ferrary[29][12] = 9'b100000100;
assign ferrary[29][13] = 9'b101001000;
assign ferrary[29][14] = 9'b101000100;
assign ferrary[29][15] = 9'b100000000;
assign ferrary[29][16] = 9'b101101000;
assign ferrary[29][17] = 9'b101101101;
assign ferrary[29][18] = 9'b101001001;
assign ferrary[29][19] = 9'b100100100;
assign ferrary[30][4] = 9'b100101001;
assign ferrary[30][5] = 9'b101110010;
assign ferrary[30][6] = 9'b101101101;
assign ferrary[30][7] = 9'b100000000;
assign ferrary[30][8] = 9'b100000000;
assign ferrary[30][9] = 9'b100100100;
assign ferrary[30][10] = 9'b100000100;
assign ferrary[30][11] = 9'b100000000;
assign ferrary[30][12] = 9'b100000000;
assign ferrary[30][13] = 9'b101001000;
assign ferrary[30][14] = 9'b101000100;
assign ferrary[30][15] = 9'b100100100;
assign ferrary[30][16] = 9'b101101000;
assign ferrary[30][17] = 9'b101001000;
assign ferrary[30][18] = 9'b101001001;
assign ferrary[30][19] = 9'b100100100;
assign ferrary[31][4] = 9'b101001001;
assign ferrary[31][5] = 9'b110010010;
assign ferrary[31][6] = 9'b101101101;
assign ferrary[31][7] = 9'b100000000;
assign ferrary[31][8] = 9'b100000000;
assign ferrary[31][9] = 9'b100000000;
assign ferrary[31][10] = 9'b100000000;
assign ferrary[31][11] = 9'b100000000;
assign ferrary[31][12] = 9'b100000000;
assign ferrary[31][13] = 9'b100100100;
assign ferrary[31][14] = 9'b101101001;
assign ferrary[31][15] = 9'b101101101;
assign ferrary[31][16] = 9'b101101000;
assign ferrary[31][17] = 9'b100100100;
assign ferrary[31][18] = 9'b101001001;
assign ferrary[31][19] = 9'b101001001;
assign ferrary[32][4] = 9'b101001001;
assign ferrary[32][5] = 9'b101001001;
assign ferrary[32][6] = 9'b100100100;
assign ferrary[32][7] = 9'b100000000;
assign ferrary[32][8] = 9'b100000000;
assign ferrary[32][9] = 9'b100000000;
assign ferrary[32][10] = 9'b100000000;
assign ferrary[32][11] = 9'b100000000;
assign ferrary[32][12] = 9'b100000000;
assign ferrary[32][13] = 9'b100000000;
assign ferrary[32][14] = 9'b100100100;
assign ferrary[32][15] = 9'b101001000;
assign ferrary[32][16] = 9'b100100100;
assign ferrary[32][17] = 9'b100000000;
assign ferrary[32][18] = 9'b100100100;
assign ferrary[32][19] = 9'b101001001;
assign ferrary[33][4] = 9'b101001001;
assign ferrary[33][5] = 9'b100101001;
assign ferrary[33][6] = 9'b100000000;
assign ferrary[33][7] = 9'b100000000;
assign ferrary[33][8] = 9'b100000000;
assign ferrary[33][9] = 9'b100000000;
assign ferrary[33][10] = 9'b100000000;
assign ferrary[33][11] = 9'b100000000;
assign ferrary[33][12] = 9'b100000000;
assign ferrary[33][13] = 9'b100000000;
assign ferrary[33][14] = 9'b100000000;
assign ferrary[33][15] = 9'b100000000;
assign ferrary[33][16] = 9'b100000000;
assign ferrary[33][17] = 9'b100000000;
assign ferrary[33][18] = 9'b100100100;
assign ferrary[33][19] = 9'b101101101;
assign ferrary[34][4] = 9'b100101001;
assign ferrary[34][5] = 9'b100101001;
assign ferrary[34][6] = 9'b100000100;
assign ferrary[34][7] = 9'b100000000;
assign ferrary[34][8] = 9'b100000000;
assign ferrary[34][9] = 9'b100000000;
assign ferrary[34][10] = 9'b100000000;
assign ferrary[34][11] = 9'b100000000;
assign ferrary[34][12] = 9'b100000000;
assign ferrary[34][13] = 9'b100000000;
assign ferrary[34][14] = 9'b100000000;
assign ferrary[34][15] = 9'b100000000;
assign ferrary[34][16] = 9'b100000000;
assign ferrary[34][17] = 9'b100000100;
assign ferrary[34][18] = 9'b100100101;
assign ferrary[34][19] = 9'b101101101;
assign ferrary[35][4] = 9'b100100101;
assign ferrary[35][5] = 9'b100101001;
assign ferrary[35][6] = 9'b100100101;
assign ferrary[35][7] = 9'b100100101;
assign ferrary[35][8] = 9'b100100101;
assign ferrary[35][9] = 9'b100100101;
assign ferrary[35][10] = 9'b100100101;
assign ferrary[35][11] = 9'b100100101;
assign ferrary[35][12] = 9'b100101001;
assign ferrary[35][13] = 9'b100101001;
assign ferrary[35][14] = 9'b101001001;
assign ferrary[35][15] = 9'b100101001;
assign ferrary[35][16] = 9'b100101001;
assign ferrary[35][17] = 9'b100100101;
assign ferrary[35][18] = 9'b100101001;
assign ferrary[35][19] = 9'b101101101;
assign ferrary[36][4] = 9'b100100100;
assign ferrary[36][5] = 9'b100101001;
assign ferrary[36][6] = 9'b100101001;
assign ferrary[36][7] = 9'b100100101;
assign ferrary[36][8] = 9'b100101001;
assign ferrary[36][9] = 9'b101001001;
assign ferrary[36][10] = 9'b101001101;
assign ferrary[36][11] = 9'b101101110;
assign ferrary[36][12] = 9'b101110010;
assign ferrary[36][13] = 9'b101110010;
assign ferrary[36][14] = 9'b101101110;
assign ferrary[36][15] = 9'b101001101;
assign ferrary[36][16] = 9'b101001001;
assign ferrary[36][17] = 9'b100101001;
assign ferrary[36][18] = 9'b100101001;
assign ferrary[36][19] = 9'b101001101;
assign ferrary[37][4] = 9'b100100100;
assign ferrary[37][5] = 9'b100101001;
assign ferrary[37][6] = 9'b101001101;
assign ferrary[37][7] = 9'b100101001;
assign ferrary[37][8] = 9'b100101001;
assign ferrary[37][9] = 9'b101001001;
assign ferrary[37][10] = 9'b101001101;
assign ferrary[37][11] = 9'b101101110;
assign ferrary[37][12] = 9'b101110010;
assign ferrary[37][13] = 9'b101110010;
assign ferrary[37][14] = 9'b101110010;
assign ferrary[37][15] = 9'b101101110;
assign ferrary[37][16] = 9'b101001001;
assign ferrary[37][17] = 9'b101001101;
assign ferrary[37][18] = 9'b101001001;
assign ferrary[37][19] = 9'b101001001;
assign ferrary[38][4] = 9'b100100100;
assign ferrary[38][5] = 9'b101001101;
assign ferrary[38][6] = 9'b101101110;
assign ferrary[38][7] = 9'b101001001;
assign ferrary[38][8] = 9'b100101001;
assign ferrary[38][9] = 9'b101001001;
assign ferrary[38][10] = 9'b101001101;
assign ferrary[38][11] = 9'b101110010;
assign ferrary[38][12] = 9'b101110010;
assign ferrary[38][13] = 9'b101110010;
assign ferrary[38][14] = 9'b101110010;
assign ferrary[38][15] = 9'b101110010;
assign ferrary[38][16] = 9'b101001101;
assign ferrary[38][17] = 9'b101110010;
assign ferrary[38][18] = 9'b101001101;
assign ferrary[38][19] = 9'b101001001;
assign ferrary[39][4] = 9'b100101001;
assign ferrary[39][5] = 9'b101101110;
assign ferrary[39][6] = 9'b110010011;
assign ferrary[39][7] = 9'b101001101;
assign ferrary[39][8] = 9'b100101001;
assign ferrary[39][9] = 9'b101001001;
assign ferrary[39][10] = 9'b101001101;
assign ferrary[39][11] = 9'b101110010;
assign ferrary[39][12] = 9'b101110010;
assign ferrary[39][13] = 9'b110010011;
assign ferrary[39][14] = 9'b110010111;
assign ferrary[39][15] = 9'b110010011;
assign ferrary[39][16] = 9'b101101110;
assign ferrary[39][17] = 9'b110010111;
assign ferrary[39][18] = 9'b101101101;
assign ferrary[39][19] = 9'b101001101;
assign ferrary[40][4] = 9'b101001101;
assign ferrary[40][5] = 9'b101110010;
assign ferrary[40][6] = 9'b110010111;
assign ferrary[40][7] = 9'b101110010;
assign ferrary[40][8] = 9'b100101001;
assign ferrary[40][9] = 9'b101001001;
assign ferrary[40][10] = 9'b101001101;
assign ferrary[40][11] = 9'b101110010;
assign ferrary[40][12] = 9'b110010011;
assign ferrary[40][13] = 9'b110010111;
assign ferrary[40][14] = 9'b110111111;
assign ferrary[40][15] = 9'b110010111;
assign ferrary[40][16] = 9'b110010010;
assign ferrary[40][17] = 9'b110010011;
assign ferrary[40][18] = 9'b101110010;
assign ferrary[40][19] = 9'b110010010;
assign ferrary[41][4] = 9'b100101001;
assign ferrary[41][5] = 9'b101001101;
assign ferrary[41][6] = 9'b110010011;
assign ferrary[41][7] = 9'b110010111;
assign ferrary[41][8] = 9'b100101001;
assign ferrary[41][9] = 9'b101001001;
assign ferrary[41][10] = 9'b101001101;
assign ferrary[41][11] = 9'b101101110;
assign ferrary[41][12] = 9'b110010011;
assign ferrary[41][13] = 9'b110111111;
assign ferrary[41][14] = 9'b111111111;
assign ferrary[41][15] = 9'b110111111;
assign ferrary[41][16] = 9'b110010010;
assign ferrary[41][17] = 9'b110010010;
assign ferrary[41][18] = 9'b101110010;
assign ferrary[41][19] = 9'b101101101;
assign ferrary[42][4] = 9'b100000000;
assign ferrary[42][5] = 9'b100100101;
assign ferrary[42][6] = 9'b101110010;
assign ferrary[42][7] = 9'b110111111;
assign ferrary[42][8] = 9'b100101001;
assign ferrary[42][9] = 9'b101001101;
assign ferrary[42][10] = 9'b101001101;
assign ferrary[42][11] = 9'b101101110;
assign ferrary[42][12] = 9'b110010011;
assign ferrary[42][13] = 9'b110111111;
assign ferrary[42][14] = 9'b111111111;
assign ferrary[42][15] = 9'b111111111;
assign ferrary[42][16] = 9'b101110010;
assign ferrary[42][17] = 9'b110010010;
assign ferrary[42][18] = 9'b101101101;
assign ferrary[42][19] = 9'b100100100;
assign ferrary[43][5] = 9'b100000100;
assign ferrary[43][6] = 9'b101110001;
assign ferrary[43][7] = 9'b110010111;
assign ferrary[43][8] = 9'b101001101;
assign ferrary[43][9] = 9'b101001101;
assign ferrary[43][10] = 9'b101001101;
assign ferrary[43][11] = 9'b101110010;
assign ferrary[43][12] = 9'b110010011;
assign ferrary[43][13] = 9'b110010111;
assign ferrary[43][14] = 9'b110111111;
assign ferrary[43][15] = 9'b110011111;
assign ferrary[43][16] = 9'b101110010;
assign ferrary[43][17] = 9'b110010010;
assign ferrary[43][18] = 9'b100101001;
assign ferrary[43][19] = 9'b100000000;
assign ferrary[44][6] = 9'b101101101;
assign ferrary[44][7] = 9'b110010010;
assign ferrary[44][8] = 9'b101001101;
assign ferrary[44][9] = 9'b101001101;
assign ferrary[44][10] = 9'b101001101;
assign ferrary[44][11] = 9'b101101110;
assign ferrary[44][12] = 9'b101110010;
assign ferrary[44][13] = 9'b110010011;
assign ferrary[44][14] = 9'b110010111;
assign ferrary[44][15] = 9'b110010011;
assign ferrary[44][16] = 9'b101110010;
assign ferrary[44][17] = 9'b110010010;
assign ferrary[44][18] = 9'b100100100;
assign ferrary[45][6] = 9'b100000100;
assign ferrary[45][7] = 9'b101101101;
assign ferrary[45][8] = 9'b101001101;
assign ferrary[45][9] = 9'b101001001;
assign ferrary[45][10] = 9'b101001101;
assign ferrary[45][11] = 9'b101101101;
assign ferrary[45][12] = 9'b101101110;
assign ferrary[45][13] = 9'b101101110;
assign ferrary[45][14] = 9'b101110010;
assign ferrary[45][15] = 9'b101101110;
assign ferrary[45][16] = 9'b101101101;
assign ferrary[45][17] = 9'b101101101;
assign ferrary[46][7] = 9'b100100100;
assign ferrary[46][8] = 9'b101001001;
assign ferrary[46][9] = 9'b101001001;
assign ferrary[46][10] = 9'b101001001;
assign ferrary[46][11] = 9'b101001001;
assign ferrary[46][12] = 9'b101001101;
assign ferrary[46][13] = 9'b101001101;
assign ferrary[46][14] = 9'b101001101;
assign ferrary[46][15] = 9'b101001101;
assign ferrary[46][16] = 9'b101001001;
assign ferrary[47][8] = 9'b100000100;
assign ferrary[47][9] = 9'b100100100;
assign ferrary[47][10] = 9'b100100101;
assign ferrary[47][11] = 9'b100101001;
assign ferrary[47][12] = 9'b100101001;
assign ferrary[47][13] = 9'b100101001;
assign ferrary[47][14] = 9'b100100101;
assign ferrary[47][15] = 9'b100100100;
//Total de Lineas = 694
endmodule

