
always @ (*) 
	
	begin 
	case (~iConteo_Tiempo_Llenado)
		
		9'b000000000 : iSelect = 15'000000000000000;  // APAGADO
		9'b000000001 : iSelect = 15'011000110101110; // END
		9'b000000010 : iSelect = 15'000000000000000; // 0
		9'b000000011 : iSelect = 15'000000000000001;// 1
		9'b000000100 : iSelect = 15'000000000000010; // 2
		9'b000000101 : iSelect = 15'000000000000011; // 3
		9'b000000110 : iSelect = 15'000000000000100; // 4
		9'b000000111 : iSelect = 15'000000000000101; // 5
		9'b000001000 : iSelect = 15'000000000000110; // 6
		9'b000001001 : iSelect = 15'000000000000111; // 7
		9'b000001010 : iSelect = 15'000000000001000; // 8
		9'b000001011 : iSelect = 15'000000000001001; // 9
		9'b000001100 : iSelect = 15'000000000101010;// 10
		9'b000001101 : iSelect = 15'000000000101011;// 11
		9'b000001110 : iSelect = 15'000000000101100; // 12
		9'b000001111 : iSelect = 15'000000000101101; // 13
		9'b000010000 : iSelect = 15'000000000101110; // 14
		9'b000010001 : iSelect = 15'000000000101111; // 15
		9'b000010010 : iSelect = 15'000000000110000; // 16
		9'b000010011 : iSelect = 15'000000000110001; // 17
		9'b000010100 : iSelect = 15'000000000110010; // 18
		9'b000010101 : iSelect = 15'000000000110011; // 19
		9'b000010110 : iSelect = 15'000000001000000; // 20
		9'b000010111 : iSelect = 15'000000001000001; // 21
		9'b000011000 : iSelect = 15'000000001000010; // 22
		9'b000011001 : iSelect = 15'000000001000011; // 23
		9'b000011010 : iSelect = 15'000000001000100; // 24
		9'b000011011 : iSelect = 15'000000001000101; // 25
		9'b000011100 : iSelect = 15'000000001000110; // 26
		9'b000011101 : iSelect = 15'000000001000111; // 27
		9'b000011110 : iSelect = 15'000000001001000; // 28
		9'b000011111 : iSelect = 15'000000001001001; // 29
		9'b000100000 : iSelect = 15'000000001100000; // 30
		9'b000100001 : iSelect = 15'000000001100001;// 31
		9'b000100010 : iSelect = 15'000000001100010;// 32
		9'b000100011 : iSelect = 15'000000001100011;// 33
		9'b000100100 : iSelect = 15'000000001100100;// 34
		9'b000100101 : iSelect = 15'000000001100101;// 35
		9'b000100110 : iSelect = 15'000000001100110;// 36
		9'b000100111 : iSelect = 15'000000001100111;// 37
		9'b000101000 : iSelect = 15'000000001101000;// 38
		9'b000101001 : iSelect = 15'000000001101001;// 39
		9'b000101010 : iSelect = 15'000000010000000;// 40
		9'b000101011 : iSelect = 15'000000010000001;// 41
		9'b000101100 : iSelect = 15'000000010000010;// 42
		9'b000101101 : iSelect = 15'000000010000011;// 43
		9'b000101110 : iSelect = 15'000000010000100;// 44
		9'b000101111 : iSelect = 15'000000010000101;// 45
		9'b000110000 : iSelect = 15'000000010000110;// 46
		9'b000110001 : iSelect = 15'000000010000111;// 47
		9'b000110010 : iSelect = 15'000000010001000;// 48
		9'b000110011 : iSelect = 15'000000010001001;// 49
		9'b000110100 : iSelect = 15'000000010100000;// 50
		9'b000110101 : iSelect = 15'000000010100001;// 51
		9'b000110110 : iSelect = 15'000000010100010;// 52
		9'b000110111 : iSelect = 15'000000010100011;// 53
		9'b000111000 : iSelect = 15'000000010100100;// 54
		9'b000111001 : iSelect = 15'000000010100101;// 55
		9'b000111010 : iSelect = 15'000000010100110;// 56
		9'b000111011 : iSelect = 15'000000010100111;// 57
		9'b000111100 : iSelect = 15'000000010101000;// 58
		9'b000111101 : iSelect = 15'000000010101001;// 59
		9'b000111110 : iSelect = 15'000000011000000;// 60
		9'b000111111 : iSelect = 15'000000011000001;// 61
		9'b001000000 : iSelect = 15'000000011000010;// 62
		9'b001000001 : iSelect = 15'000000011000011;// 63
		9'b001000010 : iSelect = 15'000000011000100; // 64
		9'b001000011 : iSelect = 15'000000011000101;// 65
		9'b001000100 : iSelect = 15'000000011000110;// 66
		9'b001000101 : iSelect = 15'000000011000111;// 67
		9'b001000110 : iSelect = 15'000000011001000;// 68
		9'b001000111 : iSelect = 15'000000011001001;// 69
		9'b001001000 : iSelect = 15'000000011100000;// 70
		9'b001001001 : iSelect = 15'000000011100001;// 71
		9'b001001010 : iSelect = 15'000000011100010;// 72
		9'b001001011 : iSelect = 15'000000011100011;// 73
		9'b001001100 : iSelect = 15'000000011100100;// 74
		9'b001001101 : iSelect = 15'000000011100101;// 75
		9'b001001110 : iSelect = 15'000000011100110;// 76
		9'b001001111 : iSelect = 15'000000011100111;// 77
		9'b001010000 : iSelect = 15'000000011101000;// 78
		9'b001010001 : iSelect = 15'000000011101001;// 79
		9'b001010010 : iSelect = 15'000000100000000;// 80;
		9'b001010011 : iSelect = 15'000000100000001;// 81
		9'b001010100 : iSelect = 15'000000100000010;// 82
		9'b001010101 : iSelect = 15'000000100000011;// 83
		9'b001010110 : iSelect = 15'000000100000100;// 84
		9'b001010111 : iSelect = 15'000000100000101;// 85
		9'b001011000 : iSelect = 15'000000100000110;// 86
		9'b001011001 : iSelect = 15'000000100000111;// 87
		9'b001011010 : iSelect = 15'000000100001000;// 88
		9'b001011011 : iSelect = 15'000000100001001;// 89
		9'b001011100 : iSelect = 15'000000100100000;// 90;
		9'b001011101 : iSelect = 15'000000100100001;// 91
		9'b001011110 : iSelect = 15'000000100100010;// 92
		9'b001011111 : iSelect = 15'000000100100011;// 93
		9'b001100000 : iSelect = 15'000000100100100;// 94
		9'b001100001 : iSelect = 15'000000100100101;// 95
		9'b001100010 : iSelect = 15'000000100100110;// 96
		9'b001100011 : iSelect = 15'000000100100111;// 97
		9'b001100100 : iSelect = 15'000000100101000;// 98
		9'b001100101 : iSelect = 15'000000100101001;// 99
		9'b001100110 : iSelect = 15'000010000000000;// 100
		
	default: iSelect = 0; // Valor por defecto
	endcase // Fin del case                                                        
	
end // Fin del bloque always
